PK   ��dXqC,&'  ��    cirkitFile.json�}[�9��_1j^�*��;鷝Ng������QH)3��T��*U_���~��LI�$S!E���c�c+�F�c0��巻m�S����l������z�t�V���ն��:������~z�m���>~�{�[�w���cS�6?~�<5O��v%��h���}Y����Ԣ]	��RW�������.h�Ʈh��nh���h������;A� "O�'��D�	"�~��?Iğ��="�$��?Iğ$�O�'���D�)"�Tmh}c�-lX�
��%�X6!�fel�j�Q?�l�VF�b�Dʕ+BeUQ/�қUU���1���hx�ߠ���Ş�5(�|�A����=�eP���b�wl��/(�/I�'bv&����LѫPiS7���W�^��K�Jj[��U�3��n(�i�n)�I����$��^:W��sn`	By)`,[I��Z�ua�ֵ��R��Vt���(�$�w��ͪI0�	q��!m&����@�O�03� . !�k�@PQ*"���?Eğ"�O���D�i"�4�����D�i"���]~UyU����e��JA����jC�H�-Lҁ��+�l��QmH��a
F5)L1ľf�}�P��ľf�}���!�zC�����m��V���U�]�vzUT���3�!T2Esm.�F�&�
�(�I��f�M���^�-;�eQ-۪h��24�
���Q�i����T�*���-��[bw��ќ#�0.���W�j]��-��}]Tm%��.W+a�]�.)F�M�qtrYأʮIe'��q�r� ��RvO�3��g|nhÕ���<1���>㳣���'F���O!�O+�!�ڎ"�8��D��X��D�j2����K��%5�WR�z%��$�P�D���CQR�]%���4���29�<��)��ę�lHT$�3�3��ʴ�+�.�X*Q�/�a��Z��e([��҃�sk(ʹ@ �K�,�-B�u�A
���ի�+��ƄҜ�5`4�ʜ��"�*�� ��\�� !h�M�H��P�s�mC(�y���X�p$�	�s��MМ��(��G���7�w�	�J@�ޑ�ݹ��IRt�(v��;�@�]����p�J+Ew��#W�Һ�N��:	e, �M�%��l���V�ܚ42�CQ��Z��EuΣ ���9G�LURT�:2AKQ�C8r�%A�$�&U�̵5r�-Euv����M�߹΅��NQ��f�]�Վ��esk��J���ۉ`��v��2�j�p���(�=Eu~Ή�Gi/�*�:��\�j��ϵ�������'��v)�E�b��Y�)�E�c��Y��1������������ÂĂŒŒ��X�X�X�X�X�X�X�X�X]D1r!����HRxl�ءp�X�\�N��E��΄[$e�r�+��Y�\�j�K��a�������� b\���1f�*�61<�G5��&�ė����Y�+۶1��K�i�t(v����N�/G581<~�rT���/G581<(�����D�)��A��A��A��A��A��A��A��A��A��A�f��yP�yP�yP�yP�;S�����QlZ�3a��O�SRb?�Gq�W%0<(6<(6L;_lx|���ŶC�i�ZSf0�C���VK��5EL���V7�+g�&�٣X�-i�hyPlyPlyP�xP�x"
��]��z�2-e�q<����bס���
�y1<(v<(v�u�,+�ږ�A��A��P\ٲ$��x������(�mI	!=OD�V�yP�y|q�AqأXB[QZ*�������������S҃+����(y�qwp�ES��rw��ES��AswęE���xLx�J�qe�.oPB�a�3W2��%�&<_��a�MG)ڙLč=}����	q�Ǚ�j�R���v)b/�^���{�x�^�G���{�w~��(�����y�aO�2�����Y�]���3�R.Q���W����	�����}du~�}�t~M	}�t~�{&t�kc�h^p3�#��k��ӏ�k�؃����3��K����K�ؓ�����C�f�����`����'�����= 7�{�m~���ڼǞ@c�r1��=S6�.���]cOz1ԋ9�\�n=�]C=��Լ��c�8��-��"E�H�,R��"űH�,R��˃^�_��_�`��`�a��a�b��bɃb��yP,yP,yP,yP,yP,yP,yP,yP�xP�.�}v�.�ǖ�
}v�.�bwB�ݢK�ؙ�g��R.v%��-�1�������-1< ����n1�����v�����rT�?�� �ŗ���-1<(����n1��A��v�AS(��bŃbŃbŃbŃbŃbŃb̓b̓b̓b��X�X�X�X�X����������0M�xPlxPlxPlxPlxPlyPlyPlyPlyPlyPl��'xPlyPlyPlyP�xP�xP�xP�xP�xP�xP옖�xP�xP�xP�yP�yP�yP�yP�yP�yP�yP�V�yP�yPxPxPxPxPxPxPxPxP��\Y��Gɔ�(�%S�dJ}�L���)�Q2e?J��GɄg�4��y\�<�TW.�+�Ǖ��J�]���nѥ\�2��]�E[�g��Rxl����g��R.�n��-���=}v�.�b�F��b@xy�{y��b��ˣ��֬��-���͍=�E��c�E��nѥ\,��֬��-���%B�ݚ@�g��R.�}v�.墻C�ݢK���س[t)<�rq@���|�����ۿ�����{�����������c�j����f[7ۻ�?P��D���os]����fJ��'�(�)���f�ݷkv_�����������ж�PTSn���I�]u�Kc�}�!ρ|�>��~��B#���ʓ���j��'�fJmg��+��Yj�fIY��h��v62AN�I�(�)��f{4r�Mڏ��qk*��wդ
��zC�+�_T����3�*��e>��-cT���u8��KA./��,̐ku��΅\�#��Nm�k�����?1���a�I���$ݔ���̰9=�����LK�vђtS�Y��/lr��%���am|��������:�N�X�Ŗ�G�9^c�|ր�X:�@\A�5�5�;������
 z���Jb�n5�@���f�[@�6{�}Ѯ�>oW�f >�x�ND|��.�c�Ĭ�g�4��.I_<8~ ��+#t�$�~�*������G�jM�Ղ�5�����fx��&�jb�n5�9�V��'����j�1�_�憄��r\�^����g�����[@�N�-�&�����U�-����P3�t�	�c��uN���n�p6���2n��3[�o1c��l��S%�s`0��݁����L��`0��"n�����������ߛ�M��,�˺�>
�@�A	"�$�+"�&�"�%�;"�'�*~� �"PP!(�T
*
���CA��"QR�(ɾ��DIE��"QR�(�H�T$J*%���D5�Dd6��]y��2�'�3�/P�3��ш�?�)p+�D��.��H��3yS#U����xEE�\̀]>;/�$-��<R��y"�>7v�rb�����7�ɀIQV1��Pi����<O�G��\p�@��s�	N ��'8T��'8�h@��*���DEE��"QQ���H�T$j*5���R���H�T$j*���΂;�Z|��ٙ<�ºI̦(��&�RB?CE���ؐ'XT*�ņ�O՟Z�?����a'��6A��<Җ������9)�fs0�#�T�[*�-㎊qG��ۺ)�%)�Ku���|����L���Qq�!�$%Ʃ��T���/��� O�<�>��EY���i���T��8�BR���*N���^��
�@N �3�BIu��w�h�i��
���b4	T@�_�I ���dL2��Ș�g�詬��/H	dL��AJ c����KJ����e&&B?v&.7�c_;��A�ς��ˤ(�����P���/�������&��o�ep�~=��)�����QJ7��o�Q��*��a�������ɣt�XS!����̊�m�3y�5�#cg�h��a��ٱ3q9_�}�̸\c`";�k�dg�2M�~��L\���o���˴,���3q�}��eg�2n�|ٙ��WA�cv&.La4����B�lv&.��'���e��~���2:�ѳ� �~�<+A\"˸�hg�2��������Ŭ�xt	�?ǳK�=�wo��h���5]d��X�ةb?�]?��sx���K�N;ݹ��v����������X��ݨ݅]|�-2r�ȡⅹw����j>��3'r�ȡ"��*r�ȡ"��:r�ȡ�D9t�БCG9L�0��D9LW��a"��&r��a#��6r��a#���)r��a#��.r���"��.r��Ẫ�.r���#��>r���#��>r��5"��!r��"G�!r��"G��k�}vM��@�s���!�^.��)�ɡ��t��]�n�"���x� �#`�=� أ`���LʏP��E̓G����#�.ǌc#q��H`��/&L0a���:���7_�����=�S�����A�d`{��뛎k�/�MGi�5�G���<��;�)ZښW�{��,6-���x�'eEnR�k��y�k:q$XC~�k:�$XC~�k:�O[�:oSM�3֐���.��!�`5��g��<j5]� XC~�j��B�����t� m�뼆5]�!XC~ k�6C���f�t�`��i�.c�k��5����>�5M���y����	>�1�'��ٓ��:�tM�Cs�wMs_s�oyMS{s��{M3�s�/~M�s�7_)v�/���j�<Ƶ���W������ҟ}R�'5���Oz������S�*��D�IL>��KL�ā-�7�LL�&���i��P61-�
'���R��7;��on�����[���79ԋ�֋�EN�EZ<��C�E(�"LKP%��
��h9m9������@N�@��i�P 9-�J �~S=>>,�MU/7�6>��n�ϻ�*_�ˡ�>������ߺ���n>6�ݺ�4?~|���5(}�m�O� ����������Ǘ����$���iJ��o�6?���{�������l��~^/��o��?^�ۦ�{�۾4P�����Z�^����d'���c�L��y^����
��{!�B��c�>��� ߝT���RΘ���骨J	�o��g��r)���{�}�������zZ��2d�w���T{�^>F�������6ra�-����>�-�)�rtrFF��t�#�"G���"�����/�a)q��#%*��h��X�WB[Z��B��7%TׄA�|tv�"Kh��r�z���"椔3%�ޞ�(G��t�}T�v�QNᘣ��1C� d�r����9�)&S��(TG���<�����w�ww�����?���û��ww��E�F@i
)K�此)|S�ES[�]U�V�}�����g���7{^�\��Y�0^�`�-�8/5L�o;ި��O)YWje#um�BὭ
�Y��-]�|�<}|ٝ0��n�jP�Zb*`��Ҵ�FV������ߚ(�/P'��X�?|X?֧f��hk�Ų�M���*��d�BX��ri�A����v��}��y:�"EPPt(Rٚ~�E��R����k�JH����9�Ư�fe�~��qJ���;�X��U�i�����_>VOu�� ��w��>�)���S'���m�����Ӧc>%�뀒�/�m����m����t/�4����I�k��E� �����V�B�hw�A�H%Ī�mr [(�lE��x�^�S�U%ji�U
`�ڕ���X�6�z�U-u���U-C� ��
fSnU�pl �Ъ���5P�]�l��绻�6���s�{�������޽{z������{���e���&R���l��7�͛��ӛ,o���i�����&-��j���m>6ծ�=�����Y�:�tV�/������ƹ�w� m���x<���H�\�߽���!��� �D,<}��'g�g���nwBۘ�ѪPK�a�����nmMp�Z��ը���ƱK�����*?�^	��J#�2�R��`z�ٔ!�����V/��ڄCs�>��p�3p����W"��f�Yذ����~o��g߽^(k����!,	`_?,���\�M��6����Z� E9��S��_�δ^���b\�e�"}���=��$����0��C-A4�A���(ݓI釆��^ɴ�}{*���qu/|�SI�U��CI�8��I��s�3$�&�RJ�����ڴ�HfD��j3I�	��N�*�](gGf!"<��t�&�RZ-�+� )�] ��:�V�"K�pY�HJk�Z;2(� �'�&��H� r�1e��J?"�yG��".����2� K}��� �4��� |WN�y�G>*v��%����	ٙo!��&M��J��+���QT_O��d��Fݫ��^NM��E�Dݱ��8������G��@]�Z��?��8�8+��t&Cg;y��'a�w��NJ%)]�j}�J�E	-ޣ�f蠸&ءy`�N���:/U��u������9����0t��0Q�G�Qu�X�= l!��ݪ���� ���.�ٷ�)A�����a��0"t�:�ʃԜ�aR��h3!��X]FsGhab5��6�9A��,�BZeT�b�J*��6Ch#EFq�0�X�M{UZqGg�!��L�MХԪ2zf��1Mi�d1�3�l3Zt)���f��.�`$ӦS��.ab�V��ɤ�6zvZi�.��ۅ�Zn���Z;2�Sa��S�$�J����8B#	��.�[��3��%�
�Z)>6��#�o%tF�.���;ѳf�vdѯ��ej8A���	��gʹ�.@|�ӝ��,����J��AKZiGä8��:�K��0���zm�j#��A̗uB�R*s�����'2J�t0���(��%����C_5q�	í:N�;"#��a>�J���}��oBh;�S��6Tr��0L���4
3b0��='�W#���8����5�,��4���ar�;A��a�ބ�*���a�|R�q2^h��e�`�:��*U.ͱ�c�M��#��a@���ިpP�*X���f/D]ڦ��#���Y���B��zj�h{*���J���:�z� ��DA����8�)aa�^����[��J�nc�O��U�}Y��|�T�D(w"ח&���P��+k����T�V�l���*_׺����ʋ��ە*��U;�-Ī�u]�ɔ���?�:�����.=��}���~�|���1B�Q�A�3{X��?
��	��/������ܟ��������Ynv�x��-����<�3�w�N�S ��YU�*�qUU�̥.�m��7�8y�6���:�y���v,�yZ� 20Ŋ�L��:���,�k�t�����0�J��`�ҭ2�~s"Nu������� ��`-�C`��U�A|=̈�dV��T�Yn�D��pG��b]	)�a�	�^@�{��`��1�.�q�>M'�4?�W�*,C�#zy���:�E��N�L'E��I�_��~B!�"�5�O����HO�����ZEwL^(�L�!��Զv�rU �V1�+/�Ư��Yݠz���y/�7??Mu��;��1����C�,|��l���pT��p�q���=t�v��-��n���Rk[��_��M��Ƃ�z�(mjUUɺ��
s���g�U`fQ1އR�ny�	U�a��PBS�Ŕ�R�ʊ�$K�qH5m��� u(� b�AJt	 (�Y-�D���a§�i�m��㍿}�{���'�t����j��?�<��q��1�8�v�ހ����O����J�&n]����PUӀ+���e���"��>um�9��vx�névq�
�����U���g����+�����/n R�V���xq�W�n5�#�h�#*U��E�D��
_���rA�a��uqj(�g;�=�5��K�ƺ���5�r��"N�I١�v�{2+���s��2�_�3�9*F�j�c��}�j�Uh��ۆ��+]�F*��L�Ȳ�L+p]s	nҠ�x7D0���q��ھt���MV��a�M�#�۸�+6Ҿfu�̉����di*76���ɴ0ן�~�ML��8Y����ؼ�,����|�n��0���^w&��s�}�����w����������~_
3r�����9�c�"�j���8�ݶ��~������A���~��7�n7���F����M��v�����sx�=1���O��(�1��m�������?1��q�~�}W�>t�~{���]<��m�]��}�џ�o��=���CFX���D ��0�HU�v3,�h�j��!A��ӻ�O �1~ڶ1��ďa�OɌË��&�����F^��GD0)O!Cz7B��t#L?�4~`0kU�ď�Ï������ͻ?��u����2�Y�y�x�U?�4~�t\U��Q�����Q���7��u��gL$Eڳ��g�R�n���gJ��dU�H���;������q����lq�a��yh�n�ёdJ&=P1FД����z�/��+����a��薙��:Ib���qv*E���x.N��|^H\1��6.7$n���3.� J�=�;��L�S��������ׇ!��_
BWX�U!H�$��7P�d��Մ,�4�V�n�H�]H�����
۸����[	=D:T>�2C&o�:��{Buz#A���`P�91�w�+����a�65N��`hL��!���h��;�`��㒐�"��66h�x�s�g�N�sD� �#�"	�hJ�FP/`�N�p�03"��t�ml27-
���Y���t:Y1�\0D쌎ա�S��m����lF�Xf�0�K�6���d�e��("��6��8'08�^��W߶��y���I�ki2�n�����Y�+۶�,�y>��k��x۸�#o˒�v�=�Lj��*3��וH<����`,�%'0�y���ml��m�E�`�Q���dE4�`e���%6	�4z��z�޼�z��=W̔���=7͔�� ��S��+�&_��Cτ(�`�}ǡ��c��P�
�ؒ7���M�]�y�?:�d��U�%`��m+����8a����+lc��M��q'7�m4g�"�W�l�G���{�L�&3$9]�:�HW8f��F��y�4��������Ř(3l	��&�6�ǹ{��V��aW��{Iq1b�)���a�)��P�	v&->&�ឞ;ch2���4�  �08����R�W̮�0�+�}��z|q�C�I
8��D�'0�̝�	���{T��կ�:_aW��4s>o��%$�|��:2d���RX�]�E�@�$P�]��73F୻���7$<�G�N|F���2q�T�6��}r��͑�LP��1�9��	޺k�|tyF����T������*��Z�vLG����+N�\cW8�n:rr[Ǿ݇;���'d2Gǒ��.�3щ�z	� ;�@>�Ȉ�+�]c�n�ht�ý0�?�wÎ.�ER�7��f%YǕ~ƃ�k��Wǆ���@'�8^(4��>١u��T�ǫ,�d"�W�!��X�ب-�Րϕ�a�_�)�
㸰�oZW��h��J�ѡ�
�L&]���c,F`���k���
k�->��p�Z8��8�A��â�U�X2,�*{��	�y`FotE���ؼ�M��	����W@�o`�L�͌�|ǒ�`/8Y?>~����5�u��|�6"����?��/��K���͏����l?��t���PK   ��dX#d�y_  G� /   images/0700f4b8-b576-4b42-8309-cd2fa5470453.pngt�8\]6,�D%M�!Z�n��wA���0ZD�G����h�(��(CB����������7Ϲf�����ګ��^k���&Ox��.����~3�m�}xr:�s�]JQ�6p�޶z������;M����g;m�!9D� ��l��t{��B9��-_���pv�IǊR��<�Q�y�㕱����y/�,�e�c���	�8��?���9v�HkG��jd+���-Ɇ1��4̦Hk�;�QVm�vPMT-/q���k�xv�Y�2��a�X���x�c}v�m.����o��#vf:�YuYS}�|V����/1��/�&⋖���G�Q������y_
QS|]�����Hp6Ƒ�&w(��m��@~�E�>d$B��O�;��ۍ���?��5�銫�r!��ߙ6]�����W,�M��p�/I?������+���3�/QW�q���6�B|8d�8$r�o��8�/�;wG�CN\I����]�v��'����!��~��j�O'�r�DOg"9��nj	=���Y���#4@�{���f���̪Qs���9��͸��8�ˊ�H��V��Pbɣ��ۖ�ER�"����g\��`�ob�-��p����q�"�C���X�[/����(����0���1� ��3����m��Iݝw��-��)����X}����}F����U0�o҈ïg�~��㹤�K�����Ò���m�X"l����޼���2J~w�����e�O��㶿��48���f5��x�C��*̪���v�e��ZZO�����WaV�y�z^�_v�����l��\aV*1"��H�o������h�aٿm�R2�� �j^#����w��k��;���YZ�]�/�ֿeI�-����d�Z��(�_̏���/���/��M��w�3<�����O�uwп,i��]�N��Ћ���M�l5����o~����-�9r��"\�_������Y!zg�K��o#���0�c�A�d��-�g���T��>����B�>5��a�xoV��� j~˒���� ���Y��Ec5�����e(����كF:Ї�o�{�	bq����8n�O�1�,p�V�E}�U��|˯�K�꥽����>ZM���MI����KE�����y���d�Maסrƥ9�x>�M#���\��WTe��@�ekS�a/R��׈������	zv��#ްt���6}f�r��a�@��`y8��O��Xa����N婔�߭"ϟy�)Ͷw�/����"�mΝ�Y^�L �f��?���O���B�����Κ��<��}�����>d9nl����2��U�]`q��#Bw�[Z��������(ڝ?��~mЅ�yE��+��F�`��_�Wߴ�dlpf��^����.����7+</}�4�E���?�*��X��R��^�>~��4�7�.p�K:�Q?�8Uݘɦ���C�䝊܏b��.�BS��M�H?��=�M+��Y�Z/;�ΎA'S����RCh��xk�> ��W����ga���I�M�X�4��Sq?���N��b	�%�s��(f�[g��8eH����}�+V7mTh�й�>j]�7��<7=���9����3C��u������eO��<m����)��(Z$���X���8��9���nw� �5�a�V�a��g���J_�鷖��&��(��kh�����م���+�u�K4�Jz���D��-�	�����= �*�N�dGCJ(s�!ˆ�S�Խ���� ��ӄf����^�@�7l�)�8
M��ӕ��*�x����I���Y�q�Ϗ����%�?��DO��A���	1��5�c�nj%k2zt ����~1=�8���������#4� �׿E?s�@U�;��G�E�~I�v� ���]��p#�n�?hCr?���fK��#O�=	� Ϫ��D��˼m��g�����~;�;Y�5��1U^��v��掄m϶jcK������~e3V�@��������z��9����!�kh�re�?Ohż�h�q���7[��@a"�d��������EQ?�]o>Wr������,{��9>G���oV۫0_��+TxT��3�=��EZ�������؎!�c;]�cQ��c������>�[3w����0U߰���\9�A�?�kJ�'ُ�!9R�xZ�f�.;���~G�M�h��2���^f�s��z~�_�����F��g��)oeR�%������w�,�s��/Q"8} ߭KH�E(U>�2\�8o��J�,�8�Ί��ü�RW��0(&;Q�]ǥ3;��8D�g9���#�<��]u]2�"�]C�Ҙ�J�.�e�,��+�����s���X�P{���v	>`��o�^�`��W��,�x��h&����ZS6��@�����h�3�q��*�W��'}�3X�+��j��[���wg�n�7Šˮ���5l�����u/C�Fɯ�ދ��]�{]v�a��Ś��y��k8�=�v�C�H%9V����Nm�Mޥ�Xb���=]�B�I$�D�7�1�k�S�hc�5ɯM�;U"t0(0f�<�+����D V9t37zJ����^
�V1�l���g�(��վ����`d
�#9oW[�1@�-�8a9�b�I�j�K���N��H7�����R�$���JL~7ʡo���{�2ɧ-���x�A��2�2J#�N^[J� ����˽�u�6���u�qK[u�"x�7r����m�
�_�ѓ��lG��҇#8��"���G�&�mٵ�d�R���FUy3�Z5^���������cjx|؞T|Q��)�_|[�S�7	nQ��\���D�:|�6Q��N�I@#��XI.�ٿ�v�_mz��5�V�^B(�t⻉���/�C�(�!���
��f���y/nj�>�:�^[�I$�+�Pu��2���h��roD���o �j(H�Ҍkp�(JĦ/���z�9��ё��U�	�VAS����5�eY��~ħ-/M� �".j�G�%􇶿%��)����<���wW3$��R��l̸�f��ط������&)M�p�t�gZ�G�o�/�j��[�4�1�g�F����#H�~ٱ�sN�}�,}��E�M}�EC�k��q����9/SP�ˡ�d�D�ifd�AMV���#�1!q�i���Z �Į�d��as�4;;���`����<\C�ltH���i�M���h�=�BꝃSH�>��3�n{϶B�|gE��/bA�Out�ܛi0�T���@�^r �
v#G�
v�eY��,C�w�_�^�u�L_o �}ۦ@Ho�c��A"��v�2��ME��.�������Fs��yٓ�����`�a�H��T��v*w[�IJ��T>%�� :#x%����rX���`*Y�`�Q�`Q����u�er�J�
��״%�F#����:���YD�eG
o��A	��c/�d����Z%�Cy����?��wh�逝p����������5���GQ���ȋ���Ė�u��I�Z$Ȕ(*�7>t����е���(`�Rf�iA���8u6�7�g�Se�q�-��G4�٨�eMjW�G���R�M(V���t����BX���-m-���'�ͷ�̑���|�y��7��}��6J )j*��[�U6k��l�����D#7`��1u)׃uF��,]t�/1\����ٗ?2�2^��*e��47�\i���S^M�g���R҉��Ϙd��e�g�y�`I&G1��Ư����O�����L�䬊�"?�vW-. g3rt�PU��7�Fz�X�|)Ү= �hl�I6HN��o&~�|a��k������1��t@٨[��(4����O�)��3��j|:�_�Je�Ha�-'bD�Xj�ȑ}";�s[zC�},�T�JE��Z���UN�z��x@�X�H�������/�/;X`�߀11��gጞ�O�5��)�&�-BGq��ӮS��/�4��~�&�w�
��a�N�9�!��Pt�v`/��z������v=1�/��G��T~Q,�nt�
Y��7��439�P��Hfj)I�y�ܑ�8���U�еN �a R�yr~�1��.����|��V��e�u��g./�D=�wf�_Lh�Y癄�K�<>eKX�t,�(�(cҡ@NTX�;<��s}�|�G��k����%PŮ~����욝WOy��R�M{]�7��s߰���U-�u(�x����4n��t�~��I�S�̞m�Z�-�=4ʳɨ�
��L����9�6�� �<K�j��a�qM�����={�p�+�I���]x�W��L]@6ؑ�'�4���TT�Ų���U��ۙ��&矇�UNrMSnL�T�]	�X�ã9�#��#�0�y&N��4fΣz#�*�߶!V����ٯi&��m\�D�~;e8}�����!&b�iZ�20��XV�c�̶p��;����v�"�;[ن�?uf��k**H��&׷C��ulL�sM&����n���E!����?�|_,G�f�DC鐷�"���������{� e����\�r 	���'嘋ݫI�䳨�=:���IIA���% �í����S�������p�q,רĦ7���n��D$���S;;F��H���vhB��P���Wǻ̀�Q��v�7|N2�Ԇ�><�m�1C1��z�)췁th�Xo<�1��.���x�J��k��G��,ȍ������9qg�g���\��vOC�q�oYP�k��v0<'��pa;��wfT	W���An#���B���0����t;�&��4h�D#[t�Y8���4�"��l3���5�T+='w��%�ɕ�����X%�Dq�@�(._�F� ���(����7�/Lc���3���fH��s�/tpP���uT�s�$��!y��\��� ����Pl�W�R�̮��Ey|��iV������W�ͷ�n�hЉҀ95
\�˳;���+�x����N�{0.��s��h���n�Q��,z�o������J�m��FrPz��  Ja���� s<��]^�5v�H�w����5 �~ϔ�ѻ�y�S������W�7e=�g�%���L��}���%Fy1\� ��C���H�3���bR���g��Y�e-&��pT�}��`���|�Ez"ø\�O�Ո���[	����=��R�L$�}r<���d�����Ƅ.�z��k�SE]�_~��%7kZ�h�C�D=񳙜�� ����z�lg��M��6��3���]�*��!Z Ky��Խ2��I&1��6���UR�99=��
"��4pu�v���(�M��ͨ� ��J}f~���4'K�Vӌnʉ���JR�/��^�Y���y���Fj7#�>DVbܴ��}|�C���V#h���ն������w^��ooP:�Gzմ�_$ϐ8��`��|���	�;�-���j����}�ElR"�^6�{*Yo��wq˫�+	�rZߵ�3$vp";6��k��O�p7AF�ۗ�/t#���_�~2y1��%�i~Ŧ$�5�=T����v3z�*�D�4���|�vY��p���"}}Oƺ�^�_���c�1'[�k�a ��F	/��27�B�=����������@,Wʘz�5��"�Ɋ�����=�
w��@U�'�s|O4���l��CI�Su��n�9j4�G=�_�+�3���Y ݌��l��)A*�����M{��f,��~&&���J�	i���jjӊ���^o�_�@#�޷L�Tn��,���kk���k��]��\4��z��(�c���� ��wV伟{8���us���
b����:oW���%���_� 6��{��Bpb�����X�G|�����ꪝh>f0]�,�A���#q�~(��!���L	MY�o��[M�)y\L�2��4k�o���f�O�z�o�E\?���%Zs�!`��w�E%u���:�qbe?G�܈o<�*�)�G��~��	�����<ςi����̀��	�颕Y�Dݴ�G.&����N���/� �WF����Q�)1�g�-(���VZ��al�!�V���u66��$t|:4O
J$�\�d��.�`�G������Y�E:��k����3�9tO'���}�2Ώ�>&��Y5�w���0�ݘ(]g�W���F� �u�{�^,�	 �nB��d��o��w!��jjar��EB�d��uy������M6��<�+��=gj��Z�'��֩�n­4�ڞuTo��۵�&��lo�W�|�<����> i̶��q��;�d^�qK*����mox�X�L]Ep�!V���Rp���>������܁����P2���5�1�C��k8B#&�S�W�K��p=5�46'�+JƸ�jg0��G�K�y����W�h����NG2�nl}?N�ѓ�ʕ�T&�!�bO��N��͊(��#N,q��H~3W<��2��KDP�W���|�&E�t��82��&P���p��X�]�/t���$~
A�0e��#hkjf+^|�Pop]���<:.�K5Gc\;���f� �G�+�My���v#{Bu����t���T8#�`[��m�M�r�϶��6sE�v�>5W��:��[|HF���Q����	�e$��y��wB��[tD�ʱ���,d���e(�m=Y�E�`����z75��	8I�v����}���k���Bř(
hq$�������Ժ�k���3D5�.F�
�P�`�`�,���!���UUT�?ol_��v�h��� �䠐������㯈��-p��?�ؘ݄~<х����c�K�_2�MJ��#�8��[��]��>9�������ù�˦חѭ�(�b���¥��׿.�p��������&��9
<�]/���t�i��E�}ߓB^�Q�YF�\�v�`[�`N��/�e8A�/��S��C7a��6�/�I%?˟�+JL�f�9J8l�g0Xu?�����1���n���VZA�;����i�i����`�]mC,3��@���Qa_'��&N5x_Ğ�;Q�o����L�~�ݣ[�;�;���KѸ�+�G�_��x��]N��bxce@K�S���_y�n�9������͘���A�8�����w����,
Co�#�?�%t��0YF!W�Q�$�x��Ȍ��pAS+O�@bE�~p���'���%�(�P�����#7~�Z�*՛�=���r��w�)zDNOH\���90$L+(�Ѻ�͂���
��<��a�I�%��8�[�Pgf�Ϙ�暝��g��gXeN.x��#��vk��O}�M:�j��)�4�e�m��CD�՘Z�$_�7�DX?z����l@H���u�d�����d~PB��zv�41A�I��:jo飕Yš�����R|"���z[Y~`r0���K��I��c��I||��qD>л�&��*��;���5��|��D�7X4��>ܳ�č��:���l�bp�+"���)�� �?D6�<\��Օ������o�i�K�z��ŝ�=�V6�G��1����i�sq@��FT�a/2�Y���(�~g1%l~���v�bc�������`a�b�Piu�h�x�5^�9;"1H�,}����D̕�l��So>�Y�iA�F����x$W�d|��R��oD���[kY_<�Tan�Q�j�^�t�G�kMH=��9�d&�{�N�\�z���X(4gA���%Ѥ��ع��s����X�'��&p{�N��g�s�wJi����S4�!u���M=�s ��ъ��~5"{'��d���M�5�=ɤ!�U/���n�w��aڕ� ܤ���E�Z�L9^�Va������E,f�_�.�6�v5�]��l<Zr��1�Q$��uY�w�.�w&L�'����\��٤0��hh�����@e�8�8�����G�h)�ը8�B}�^�dO!�Wu���gF�C��){4r�q�����?hJaΨΧU?��O?��Z+Q����"�0M���������=�c��F���rӌ��'Ζ3������ɬkC��N��2k�F�N�
|菨S�[��ٽ	r?Q�u��mW"��Q��E�-r�� �{�-��� ��|�(����}�W��ѣ�U�z����|�1��'������)��&�g��)z��v��Y����*rP��l���w�nwi/~����s�U��Ĕ'��&zE}�Tٞ3�*����yg����>����?ǪM}�l��Wҩ�S6=:S��ԑ�,yS��$�R}�lc�F���e�;O�B����]9��Z0p5zjm��L9�a���vM��T�;�՞���4�G��{��i�~v/ۜ��?��T��d�u����!�SUlqB!��O؍�H�Ú��I'�C���z���MƬ��u�]b��r޻{V9w@_,�#�0�]4����Q���q��S:����~���5�Y{����A�	���Q��{˂}x���I!p샹��GS9l����"��0E!G��6Y����	~w�,P��x��(�1�9���K�+��̛�e�Bs��m~{���L'E���i�����kgujN_D���l^��U��c�
]��`3���i���,��1?�%4���z�����,;�	P����c�K����rN��;�r�E���/t�c.��A�}�&�ފn�V,Xx��"�����}Iyے�>��4�B�9��~B�i�^6�����v} �(�(po��v-�>��{�d�Nf��ahB ��^=`����w1jy[d�1�zR�(��(t������]��+&�^?K�dM����g5r��ŉW凋�S�k��O6K�"!Uś������I3y��Ǽ�����C���<aƠ�޵�v�:�dOM���T0�j��s�f�0���oJ�G�����̽�T�ƽ�M@����j��/p7.�14����$ۨ���Ki>�P��L]�-������&���O'�}Y��<[�C���`�g����DRQs~�W;��$]�x�l���c�\-�����d���n@���I(D��!3�*����2=�m�QH|ፏʁCK:�u��d��+��o����"�<u
VP�]+��-�m'��S����
�'u�yI�F�����a>�BO"��3Ӣɨ-9���s�cmnF�p�� �W�-����)����F�h�&\m
R\��8����������q͑���>���{�I���Q�\�|�C	�29v\ �����I	�}3��v.. o���p�{߾��y�&
D�/��~G����}���៝�x t������e&�؈a)������U�ԓM�D�5H��t� �Xv������� �5��,�{<���C$Rf+}����]o4����ㄬ��D��}cj1��Q�gb����+�#e(�G3;_�ܫ�̱��
�� �ݧi����Y'}�c�'udY���a����Ո�c��׿X����Q1E҄�?�'R�7�?h�kh��ns3w��Lh��# ���ˍFوp�N��6qC�";ޢf�Qu��E��QqXL~W����&����?�����L�_H� �������6f�t
�\�p���'G}��W$�V7e�C��f��;�F�
�Y�Ey/�N��a���b�Į���-B٥=�7���^�!(�ZPwZZοđd�� BU�=�a�ǣK����qo:��\t�lX�\�L�֬�ݥ�PPl~��x;@����0:	0�ڋ�M���/�h4mr	���7��,z+�4٣Q��f�D��Q�c"�?jlE&�|���"��r2����s��Q�N�/?ER���K�d���i�xx����XVt�9����ޙ�h�p86�`q��?��`S�	I��e����hA�|^@UWZ~�)&p�f��
�+��f�C�c�1P~�M�d�m�x��z���r���)Wd>H0�X���s������Jt�	�S�_wBV���q���¬�c7�QKWy^�n� ��&���:G������F��Onc,@�AI$�wF���q��6�@3���P�m�{A$?����`V&�yMqn�Jh(��@U�<����z2��7(��1h~$ռڍ<�b��N>�����*¢���
���M_���lrNnGWn��:4�y������#�����`�<����HƯx��O��V�j���=�f9�H�Fw������
v�ڮ)�.��V��i��a�x�.��{,ۭ���D�m*���v�Mf�+	�V��pU3�j���"�8_�uHM�%��k�]oӓ�:K�]l��pօ6�s�{�2�&��{�̎��!�؋���;Y��o:��w�4��w�x-g�?����}�K��u�l-�"�#����E5���u�ӡ�g߉9If'���f�G��L��^����~��q{k�#�3D_F�����)��d��4�'�x��]{̷G7\��.َ'/����imB#������G��pV��ik�F!��G�H"(����xM�lk`.����t�	�u���PC6P���#�F�?!�LS$+�<����������g�S�K����˵G��s-���w.Tٯ: �Y���;"����`�1Q	膷k(N�F�ܽ{^�/k�z��_��_D��@�u�ڷ+9�����~�}n��3�a���C��W��`B�^����	~�j��M�ʋw]��{��P�}SI�غ ��p0f. ��o��\DB�،7�_S�e�1H�Y��([�cY�sZ���xD2u�|eJ\?�g��DQm�2�nKi�D��!�Fs�V�[=}���P�a�i�渧|����!OAP�UE�*p$E�л��lړ��86R��M��`˵��1�V]�m,�h�I�J��ϫ�����?�3.�َ
4�0�~LE�Gu䈖�́n���8ǣY��U#�Ӧ�e��c�k��dJ�x�O�g$՗U�Rז�	��.h�X���pD��9�bt�l�4��Sӳ4�����um(:��c�X��mcmYpv�.�t��@{���pf=0we�K�^a������x(�J�M��9�_ɢ��|�9p�o��R|�z*zX$�)�hEv�3T�h��,���`.ձ�;/�}��P�Z��,�+�nإ3�և��N�_�6 ��KDRm�g������H��<]�I�C��W�m-D7���q��5��獎�٭�����7m�5��u~���H��Y�ns��m$Ĺ^�H��lx�*��,�F����	Y:'d�Ͼ��Ҩ���8
�yg�I���; �\F��F����<g�N�U^���ƨZv���W��4��I�s�o�U>tг3K`�$� ��Z���������Z3�|��V�b�-�I��>/����3:w�!��Nj3����-=�t|���G�oxK��,-"�{t��N#t\�ڲ��~vqG�_gK��2����lz��9e��0�b2�$��ٛP�$���2�@%�� �<�Z�-�s�֡�u.5 �M�C U���1U������dܟ�����p?�f����R�{SES�=�^Oqg����)�U����3h�)L�-��	�6���� �����GT^������wBx��6����zΝ5ʒ;zYXO0��hZ���PW�ѝ�a� ��C�NR>Tpl���o�{�ץU��!^�V���e�2�]� �=�����[��I�������`oM�H���6fU�h>�5��k���Yl�5� ]k�1/S�M��1/O+s��+Ὺ��3~m�_=��(��f���3�A����o��HK��3�G�t�褎�gh�sTc�gT#0d�z��`1|�	�����w��U���h4q�M�ሰ$UT*̬(M��y�����t��G7k|�������:RN��P���ȟ�̢���Ăvv\<H����ZT����"�H�w���Л������5;�Ϻ��OU75kaF��f�x�WL?֎DAu���d��\uT5i�Q�L���U;���<Q58�"��`�q�sG{�OJ	��l�����y�5wL����O�
DN'N�҄�p	1Y�^��c`dmK{#�㵍F��Ѵ��✺>�M�R_E6G��}��iO�*&��&~�G^����b9E_�1k������ ����hܛX�g����/�P�f~�}�'��z��vy�g���Y?p����t������!&3��K�y�i�/��U3Q�^-�����6�#��Ta �͋ ۭR�h�?s���<�z�|�!O*�oh8~&C�I��#!�U���ˈ���Aw�3ϳ������)��ailI<{zH��/�,"9��MM�Wmݍx�+;�.!�b�=��G�������D���JT�Qq��z�r�Z�Q,b�z�dh,���u7�V��R�����z�1����&�5�u�aN���z<!.�<�OT�ʌ{W�����,!!!-#crh(Ҿ!�"*��Xn�^2��|���T����a�P�N���	O����I𡵵57w�Ɔ���P	��˱�Ig���%q�l��ʉ��!(��S��{�Dm%�Cӡ�![�(J��ȅJ~ʨ�.����Rl�Uʐ0���<�sfK����#6��􈊊*Ճ�a�������5���0p^�:<�q�Jxs:JN���2-5999�؇�P�T8��*�ٖҪ�s+��\��vS.?7,쎪�*��)�ıJ��3�q����Du�8�~�211����W��M�� ��͚��s���C����R�߉*�����|E��,({~�%�?�_�p�M�K�(Բ����G��~S�����%����K�i{~Ԧ��9\�*����JM8��0FŦ����>{����  ����D,�E8���Ҫ"i�{'-��0���������k�=�a���-b9�}��nT�D�����R��f���-}�?Aɝ71����PjZ��������]�h=���~�Nb5a�A4�Njǒ�Nɹz�fu������ϸ:������~0'n�N��,�W��m甄��8��J��`�bo�����f�:q;U&��ݙ�T���ro���~�����\��K�B/=�P줣��{������J��Rw҉,���RG�����)b���6],^�wÿk͏�߄�^�\�-�j`
��uhH		�l}�VUSq�`�Р���n���B�Hb�=�N���b�j�-�pdx��dwו����i0r�$ݟ��*Qkhhx��TB4L�h/�6��[r�t���GW�,�����#����MML���sg�~���̯��TL.�077-���zIQ1)��Xu!!͛MJMM6�ς�9ڣ��0�4jp���d�*��-ޚz(�pdd�Ǌl�����U/B��m�K[[���f�˗�EEE$�Ǣ��Oϲ�:^���!f=��5�եvT�5�0�{�U�$��J�| �= �8��kh�Y��?Ɓ-��ΜQ�9��Z������^��e({���5�Er;[�Rڇ5�>�g.�E���'-gZǁ��+**0L��3��Z4?1�J�a<f;[5UW�-�Ѓo�#�)()'~�����,߾���Q�
e��d՛]\��(����1�T�UM�MC�#���9@��[(���	6�:�0��4�+A�~ѥ��k��>dAf�S���aQ�Ǒ鐧�}��ԏ��h���nv�tz����WMb[l� ��b���
u�ݼ��8��� -)�Rg&}��s�s�f�f��kcS̚4�*��\9�)Z�&q�1:�"zD�����61 7��}��<�D}���V�#�.u[��5 ���7�:.+w�;~	Ϛ�G��-��\��n�zP�aR�(�Ϋ��_�˔�
~��@�Մ9/*��}j@�cʸ&�%��|�/}�@xB{�����Ǐ�
�iH�)�3�~u�oLm�؏Z�M&���Howos���+˗��=<:*����~f�_����k�t���,%���W8�
����u��,�57�H��}ѫ�\�����$7�*�F(��N�ez߿q�R�������]���7îT�%���޻�u�E/��ә���gFI��>Њv�
�9�JQ��"?-��.���{gI�2�r�N��ۯ ����ڊ���}B[.�B���3��2�����}�k�߼1��.Ô�����-��ӝ���ѷ�r_<�X��3ӻ���=�v�{x�y�%=ۛ�/��нVf�;3�NB�A�����]LE]�H��^?�z���zn
��)Ȅ������E���g+��{.A�Q��c���J���;��d����P���E�XX4�(fb���'��9z�\=��o�p=z����/G� �WÝGf����',�0j@��v�����0xhd��2���o�L��T&�=%��ᩊ+<�=K�;K;�?���!���mU7C'�a��� ��>�3��C����0����&	�T�e�2(44T�x"%5U����r�~��k��T&�_�\��ć(��LLL%ӛ��Y��ѱJ�\bbQ&���ԑL�ڍ�:�_�^�����~7����@�9��lQ�ިB`��Z ��B �x�|�cJKK�$�W���?j�|��Jq�����].�����G~���^�:����D{�(ʯ
d_u���XN���l�(����fff4���I���em �s5���z�W]���N�gk�T��B@�&�����ր-P ��WG��C��u��Iq~�o�fq ��`�p]�L>r�\*)����	��&}!�PB�I�{Կx!�3����$V�wli{]I<�c��1+p�G5>$�bbp'ȧn���r�-�H����wr��^���]�E�������Xj�Ph)edd���P����̿\I��X
x"�T�r��j�lgpn<�5&[c�=5E�.����=푄��`�)}3(&����M\�E�T���!X�p������"7��s�q*�I��Fe�
��&<b���f�f������V f�gq��<eԲ����aá��,�ʿGp���N9���8����i�%U�#�4��@�h*T�4�cɢM���n�wt$p7��G٤{K� y��Z���)�6�B�;����~X�GF��cb�8�|䀘���W�)���5q%�KE_�{_,����gOR���@�O^1��]���W"~�&�1���q;��b*��맽G�J���>�'V�d�R�NU��̶*����ʻOFY%/�:��Kzo|����3D���;��������Ŀ6C`�_�&�����*,�v�9���{�\�c�Ƹ�����������H��k��ø���srF��Z�;Ko9j�i���^(Lu'�w�1� �B]//���� ��ae)����x�x�g��Q�íI�����P�NR找/j�m��u�o=e�&�˨w�*ߥ�'��}��;;JK�:o��jTMI�](�G��$�t�jŢ7P&g�o��2�����6�U=,D�z��}-�	:|o%�w�3B)'�l�Ҟ���f�����vt|J�ޟ���^��❉2���9&�O)�B��'X5W�xu�(������ZJ|�����-��lğ����-���s�er�ѝ�e�����7TTI���X��#�5s�ʒX� p1���ϻ�WI����1΁���y��v�Ǘ}�eu�,o.��ޒ�q ���� 놘����0�ʄ��Q7A`�3�I]y��Di_���Z� s] ���P�(4Y���n�y-���G����,f�ӗ�_ߟ�:���e��j���U���}�ޘ�ɱ��/��/� 縺�pAxџB�#8�7�6}
����(8��m�T�y���m�[����7� $�[�� �aS>��^5�Bq��؏;#�}o���vww�x|Wuqh0R`L�
������w< ��r�h A	 ~J]y?O(�@iR(��B�D�ybs���Id����P��h10Ј3$(	�T�$�S��]����v��ڑ�������/�؅�J�ez���2�U����;�?}�0��1�^�:;;�8�w֚��`(�'����j9�\c�l}-�g��I�����{4��)��H([��,���Lba�IDY8���W�xg�H���/�{n�?h�C$Q�4��!8��՛i��c����Y}��,�cr�UQg|��ʍW�'�=B�||�V4<����kHfZ�X�bC�غ�US�%?�N�&ڨ��*�[[[z�"��?1���q؉U1�z��ɸ�Ł`�����1��!�Iħ����T|~���(�;�i2�bY-RW0)��u��-z�f`����:F�����1��APse�` �Va�<���i"��~W}�:ԶL��F��Q�X��B�ź������v�nTNo6�s�3n L��*��צq�򚘆��}�W�X0������!,�w��^ ��+�c�#�_}#Z̼�2����t���'�9l�Q^�&���|�`n����q��䧬�� aN|/�_^�P��jpx��뻨;�]��Eo�HK(򪢌U= ��	tGd���l@�L)
���'�}�g6vQ$E�.z�tg���Y����t0�Jʂĭ��2�w璳�}����W�7P �e:�m��+}����$7ns�a�q��=T��ë���:�}���9��c�涗��V!11j��#��M�ZK`;oV��w�L)������K��li���mm�����i��,����� d����P�gM����g~ �$rB#�l4�p��ygUrQ6/�cO�C���KDD�t�t������j��&�kax���8w?�y��������e1ʭ%r�ɹ�d��#[K�4�/�|s(�TDD�j
᎟�cu��ɏn*�`��Uܛ�����(�8y���������>Jl�}��)c皬�:��>-��Q�����W�R�>���OU��u��x�����+��~߷GJF�t	���n��R"R�Fa�4HH�t���.)A�������p<��S�}_�c�K�[י ����ڬ�K"t�V�Yw�8G��#��_�B�����[lؽ��3���a�&8(��3y�s��G�!�����[LX�va����>>� me���Z�?8w9%��c�]� ��yS��5��FKGW�~ �W��Џ��HZjh���9u��-��̒��1����eFtY!j�����(�QαM|�>l����FW�-iaƙ�v���G�y��,9�����)?~-� ����o3�2k!�}�GJ�ۖ�NK�H0i6�S�җ9�Cl�?(0�7�
j6�/�)P����5I|����< �nv��Q������|����-bՕ�Eݺܽ��C!����W4����SB�),	�ʅ��ݚk&ǌڜ(`w�K³9�ǹ�������b�YY��΋��ߴ�� ����U�EM�Y�k�7I�kN�HNZa�� ������z�4U��q8��_1!��!���x �5�ݻ&_��׻�g��Y�y�8y&W��n��E����`�۽����+� ��ŝ��o?\}V|X�ݛ=eY�ݸ��^�6��W��ݭX9 ����0���K°���R��w����^��s1*fGޚ��Ic�b�������h�+0[	�*�z.jO�����߿]|�hӪH0?v��ż�
�Y��@N�>v��X-�@$�U���Ȍ��O�'�n���-v'y��-�F�S=k�H�U����dF�g��W1n��K��?�/���iD(�%���XQ�T�c�+�1\��}g�ꞙ���ͧ5���h�C����G��W�}��y�����Z��:��y��=%�����%z�U��T.��PT֊t�a��ý�����X١����ᔬO9j��$SݣM���(7(���@Ï�:��=�s�C���g��Y]|�N!�t����V]����D._�9������Ȇ��w��6��],u��s��-�c��[���9i�;�1RLx�U��� thc��DN"b	���p'���[��{M�'/��%�"�����FO��6(O@[x,�_�']M��5+9ի�Bz~�u����|BW�W������f�s���z�P��@��'ٛ1�=�Π��?����O�p���,w}IRQ�3�󐎴���`���P�[:�%��0�CP<�psܗ���,�C8�!U�/LT���n �i�X��jd%=q�	R---��r>>�c;9�g��C$gd�TZ��LJ۸n����06�4X3�/�9¿��������G�B��OCP�ff�<���N}���|�|��z�!'+��就)�~דP��������qß�j3U_θ��&x5�NK������m���4�NR-�_�?9�j2%���l]#�k$Y5xaل{�.N	0׳��P^�t�F�42,k��֧q�?4��2J�|��{�d~8�~LP�����:��{��f�7���i7�N�c!aa���sPn����d�i�?�}�coO���ފ�G����4�no��@�p8)Ea�'GQ�l��&L\�Z�5�Ʋ��+���r��y��Z� �3�C�Px��>PC��%����c�B� ��y���E%�*
��#�T��Vqw*>--�M+_|�x�x+�
��L�_'�OMl+	��J�z�B!��,\"��G�㉺U�����v��;}���P8�ȎxM�a����&��/bM����7ް�����=��؎WΝj�lj�~j!*)�TTك���ITLL�o�ԓ��&<_OCR���/wvL*�쉾�������,����Qp�dk6�p�"޳A���/8?�M�ӾJg���N(�#�<�t]�I6����,�����VwX�[<�~��v1r_��~�!Ub�ݥm�P��V��� �8�Bݘ�������q��ߺ � ;����Mm��"x����*��lo�î���m��x���l�K5�R�څI���I([DB���є���R�,�'���?��>^b(��Wd��d��Ԁ��"`u|��K�7���!�CZ�	���~cl�\�} ���q���N����jr~�����{Q�{D�v�1�j����P��\?�����H�RX��0��g�o���w���Yq���LÌ�ˣm��V����#�H��>���?Rb��.��$p���/h���FmPྐྵp�O�<5Hw�Җ��UCgړv�lvz�J���,0��v��b��T ����2]���s��JK�ˁl��s�uFS���h�f�$e�D��k ��9�Uu��㳮-K���P��VTɶH/�--m���[<�f��Z����	:0� �=��`��e���(E��d+D(�ӑiXbF�s�o�|a�8�>,0��H�怼�:K3������ׯ����"����z��9�����^�?�zZ��̥����yT������N�*C� ��M�"4!@!�{��k\8���d��T�T�a)�ac�������*K^�'�=}_�.�w�i$�r���&�JC���lp��pp�(��Z.�פ��U�L�R �'2�\`�;�u��#��q�O�׊u,8'USQ��R����y{{�^�ʲ�'�LżǇA�]s�p��<BB��.�D��8��v�{�giפ@��8ʰ�ǅW3�z��G�*ibC�Uז�_�2m�(P�+V��J�^���(' NOb[����HUH����}�/��%76��#���ҝy��|Z_g�q'�a��q�R�}�]�i�x0rWx���mNNR�(���)EsU���9�o�
{���؁�(���X�����üz`]�Ra�,�9��:w�v�{�EB _�����fG�a���F�����75㰪B����#B���~ꑰ�Z&RDȘ3u�Fs��Bo�P9�a����L�yl+C��j#�+o��h�d���nh
h�OQVVDx8��+A\-�mw��n�~֌E��$����C�#�RII*��_~�ܞ�L�ι_�}��Sz�}﹢�r�|!y�v�}�Y�(��z��,�巛m�V�@�R�Xf��ϟ�.7��TA���ȍ�͛�@��Sv�Z����3�i�v[1���ܹ�HH�O�x?�������FO-s�������b��?�-;yX�����1
�c@s��<t$aĜ����q��QbC{�$�u��A������:��rs��<o�ExHftA����5��AhWe����:�CM�:Ô�]7GX�c�m�A��vĕ��
���t����
Ayy���s��ۨ`#��n� ҪD��*@��5wh�j{����ب�� ��!�w��)��e�<H���f.�t�{IO�= ��Jy��mW;�̿���j]GP����{zO/#, \���0�O����P)}��.��m9���LU���=lR��t2]_FD��M>flC��C��}X��"�_�|��UP%ɷ������3hJ������bqף�4���b�
��?ym���ˑui<&6C���2��־��%X8�-���cPa{���
�yA��N�~2�H��������'(u~�+خ|��c��X���8嶇�@�S68�t{O�@v��m�\8#�����z�e����E�fQ�P��G�֎R�6�����~ɪk!`�*/�}�pf�u
h�b�"ӷ��_-Guo��t�E�=5aO/z���u�l�X7H�_,^������Ҍ}�~&����p������M�e�$��)%@P��h`�58(�:k���׈�"q�Z���K3eq��{7N��i�ן�uT��?m�RN^���}���R��4�&��9�ܤ����3eg<3�A�(����i����+��5�xr���X��)W{Gy�'º�������6����Dk�{s��D�m
��#E|{������R!8 EOf~�,��iD�8ɥ^�Iq�I+�~���(�_�+�9"֤�]T\�g�*��<G��&�12c{��--Q����9�R}�Lɱ8<G׈�N��Ae}ٜ�LA���b@������
�[�Y������q��Ԣ�	�C���g�S�`�^ȯ�����sT�AS��P�p����E��W_����pa?y�?J�Eۆ�~���*��LkM����),��5^0{Ҟ�Ff;�plH3G���7�}zP�>_�5���c~�Q��2�I��R\Gj͇jX�Ȉ�e�Z��
:��8�ߍ��8*��d%��V�-8�
����������ol85h������Z��K4T㥈C}	�i^�UQ,��_���dx��x��"�W7�1��)�x:���j�Q���#n���	������¡7��QP���;h���;ſ�ۆ��zQ�#e��C�2�u��_�T��/��lb��M�~�EM��i>< ��B�
P��X�,��F5/?�ͨs��f���A3K�ѱy�p�P���c�V��x^�r�����s��U�d\{��m�������*�e�*��#���i	�U{"���:ǰ�Q��s�E�&S��:��#�[�bU�q�jT-��wHwѲI���P/#���W�Y��䄨�d4,0�"��
I�x����9
`����7���PKN�a������I/���~gV�x�S�Ιo;�?���g �XGDƖɎd(��t��U��ҺsP�M�U0Ţ�ɤ���!�<�� ���%�~�7�V R �sVF�AY��	$��������g�p�3�y.��u�ƕ�L%j�:�&N�}��[R�͢}�8��8�_���]��U�X� /�g��&�/��d���w[�t"e����¥w�sV9��"$�����C?g �wb��N�@��r e�y����	�gM��t�c<U�����:ˁ_�lB��Z�Xg�x�S'�����Żf��׻T&����*���62@���k�}�������o/�]:9�*�i7�Ģ��%��D��u	4l2:^��Y�B�֙ң�&Rxp����W�B�9��T����~���!�{N��l��\f�	�8���C҅�6�
-iB�t��k�|1�����^nb}���-�<�D������107�~Q��K�)�l��n�H��ҕ�W����u���ʒk�(A T6�.-,<���R��k�ºȐ2��iP�|�*��_ى�y�~�Q��� �Y�([:�@ȧ�}s����s�pġ�3wt��Oި�.eZ/�Ȥ|oW#њ Ȃ�3��!e}A?�Ƅ8EPn�[��K���P��C�d� �]�θ�y������^�co��\��iD�s��t]����$��c:����p�gI9��?峧��XWJy?56ڎ���n��N.<��+H�Ƌ�)o.�
le��Å�Cs��cGdЩ� 5c(���QGƅ��XM_3��Υ��-b�#���-��}淪���uA�!?��p��l�!�:KJ^��{)[(^UR�e�\��#R�%�㠕N�2;�t���7ǅc28G��4_��.(��8��\S�H
C�Y��v���	�]�!��-Hy�>c��Bۙ���,�ͅ�U�+ߢ�"�R�v�C���b��i�P�x��_t�ߌ(�?
C�~�p�RYp0֪�̡~5��$��7���^����8T(Qf�8���ф�$4������d71z��~!;L�T�)��_��~8D	�aݥb�kvB@q�2f�e�#I�����$�òz�%qO�M&�|�� ���L��NR�_@�7���qd.��0�H_v��F<_y����~�?�(z�q��H�i�P>���q`�b�p��J%�����i��\�)F*=�Bw`�T83M�J�X�G#%D�a�(+��՘����&8n�,�,yJ�s�D��k�%�"�X���3~]�NAʁPJ=��i5�"qM/y-���H�;�ϱL��� �`R��� P�P,
�pţWh4�A����P�~���mK>��&��B'����d?��]��+-��we+���%I�S�L���j?v�5��:�l�1�&�	C��Hp^��P�v�D*v������<�c4�y���� �����E�:�9��Kv^Ig����*Xj�Y�l�-���F�v���px�z�#��������fє��m��N1^�O��r"t����N�b���!�k��I�B6(������Ru�����	#�gU�=b�)��`�95� ��KCT��got���{�l��Q�i��W����j�U#f%����\�z�h7i�Չ�H�+��?b�I�_�6>s""�<�Vl1���5�_O}E��>�0���o+E��&�؛�W]��eg��`��˛������x�.F��|���좍>�1$p���4ޗ��1���㶷x�-h�ok��Yl%!�J�����0����c�HY�_U��y,_�өi$W��-�"d55�q�����C]8�4�;Taz��X��c2���6 ���u
�w:�]��N*�/?��/���ag9���p� TN�nWux�ci�*^�	j�i�&��p�R1�P�3�ɻy�]�<�0�XB��I�cM1!�"Q־N��h<g7�D;e�8��"���F����� 1 j��86%�g��u
�>il>_�)1z�H��KB�`|z-W��4�a鼝b:��I�#��2T~�$ S��$�)xTY*�i�R�{�Q�|���wKZ���� ][�9=�\ur�u;��T��*P=k������[j�<�@s���ɑ�\�<���3SC2��.G)G�2���Y<y.�Q����㡇t$�Zy_�XF`H��F?h�bz��U��F6l�(�L����*����%rPǽ�"W��"aL<!SC�i_7ӴK6���&�ۉ�x� ��.�&�
��\�J����'���D�b*��-G5"=�p��R=�W�/Q��:����B�:�N6�D�d9���� �^��NE޳B��PD�3;Z儳�]����H�?���%� �2��v��}�vw��c��NYK�CY~%вO�p�9д1u���S�� C=L2�D�<PtQ����P$�Ԏ�~i�.��VQO����a��L鶾e�E��l����x Q-0�x?�ܭ+�^�~�x�oɬ���X�Hg�c���r�-��A�`:�6�D�pZ��0�e��^�Ԏ����qY�?6w��A��[�ѹX������D.삔
���V����j�Gb|�+�U����*;���B����X	ϷmQ���ӍI*�#�<2(���i/R��ț��Z1�y�xQ�v���hǱ�i/kJ�r��3��S���<�s��]|�g
ǫ��e�ӫ�BS��FZc���~Hr�5G�YM��3���Y�B��P�
'���A�u�yE#п�jrDx�u}��jl��:���Vp��h[�ne��f}�%=�n��|�q*��Fм�0���D��n��j�v����FћP�X/�Z�Y�Q�%?�������9��&��??��f�G[g:A�F��B`�8)�o�G�>О�J������|~>0�l�or������_�����Q�̚��k��*
H�Y;bu*�;Q�!�[w��e>� n=����(_����ɕ),=J��������$o��[�z�?�@�[~��TӁ�^���p�cM�L�G��@�,����T.�a7��r�i��6&>�@��7˅�����W���D�>Um�K	�됔Ot�Ir�Tcz��"����V{�^�)O�K
S�*����U���ؚ�V��rc7t	�8��m�f$��(0�e�})'IYL���0��R��e�)�}�LN�\�=O�$�)�eia ,9o9sV̰���s�U�Ӆ*�K�֟��m���-ƨB�҃w�`����h�Ϳ) ����:05�!\�A�IG��P6�Y�--��1캵 DC������ԏ4��A �-�I^^��e�o�2�Ϳ��WM�m��3��U��x�7�f���zӍ2Z!ԥS׆�IGl$���e
��H]fWL�!��\޲�y�"���,���O��a�@X����P�>`g?!�J��7
����T��y=hcw�KǾ~Sn�Ƀ�O� ͛y-Χ�YL%i=-ԝ/�~o8��bM�1<?ǧ��cH4V��ء9�.�W`Rf0V)kn�Je��a<�z�U1�I�� �j6;i��!�s�����TT�k�[���_t����B���f'A�/��)��ә/v<Dg�'&gCx�ke����Jȸy%Mګ޻LY�ȷQ'�8��+7 HR	w�<<�G�h����3p�L/��¹ɾ^�����H��aP����٪�ļ*h�/��n�!�����W�c-��D���T,��ZWO?��1��d��5��QȜ=��%��۾y߮J�\/���{E!���d0���P�;#�[�RA�������x�(�#t�ې�aI�n��nya�����d8�i����1+�L
���z�HL�}6e��)Mm�9n!�2"��^�C��y��PSؼlI<�<^X��$��aՄʘO����GYq�qn�ýD!�S���_ͣ7D�)�4ϣI�� �d���E��p��V�A��6����f3"�5�H:!̉���F=�|����C�5.�����w]�D�b��qpW�n~�F�dV��ϾN�c�`����G����)�#��^�n�䵝�����������@���L ۞�����a2@�]��|x����6
I0��Q�LLw���Cf���P~�Ĭb���:M�OL����:�R�`�Տt�!=�īY%N6���`�H�U����a^�$}�R�N$���'^�	n�ܼ�Σy�w@��f|ۮ?6�o�'�}��KqLǩ���:z�v��/�O�����gM>�[�vbص��\:�ߓɭ��e�U:�lw�yH�S�&��q�`���T�H��ԟS��].�\�F\���s8��J�����(i_Ix�;3CF�8:nR�}y���v�fN`�)����u>����&R�o���-��d�%�o���A�9G��[��]����F�@�n��m��T�ɺ�c���%7�a.CY� ���p��;8"��<OA��Y>��,Zt495�!������)�ـ�ۜ�s�2�s�� �7ԙ��IS{��I���^΃�S,�|�:y�lll����^�L3�943�tm�V����-i����L�(Kɲ�L���!����D�7��J����/��Y1�÷�_H��ڹ`����=ob�w(�@M�am�e�@r����޸�s�C�Ǧ���p��Uۿ��@-^� �e��E�&�e�͋���.�r�mm&Z��jQ��G�]Cm�Ь(��4����z睝���W_���﷗Yܣ�q�6��tYV�j�69�w�^+����S���B�ll��<�C3?���ٛn�Z�?x�i��~����n��p��T`NV��B�6/Y�k[Jܶ;c�,�	}H C�5���)����*g��A���=��̞G�/9V~}�SL2\s�3,�V�-����������y˱9<�GBͺ����4QC����:"8YB���;pR޶~3j��v���`�L�&2V����0�k�>���2в�m[G�+lx2Ɣ����URn{u�^�RYz�L��<ƃ��9�>h���j�� �CS���m�<"�J��ݗ	nv������D9�C�p1J:�`��qN^�	d��
�j���q%!!a�Q�U��&V�b�Ųb��DWm�F�q�����5�Mo�ɐ[�{_��L��1�[�x������8����P�Z�f�,��������h��Yf?  y�Cid�h@�]c\��Iy�m^��X7r��<����'COsg���I�i��1x�q�����0�����a-������%�M��!�#�n1?#�4�6?ELPB�]�a��`K�������^p�-�%WE.T���y�����OML�'�$V�BoaUCXrZ(�ڹ��=8�x��#>����Vs� ����t����.G��\?�����z��d�lm�2�xw=3� �{�׈���NY�&&O��;Щ<6#+�Ю�é��N*g�D.E��R����%�����S���Ȇ���:H��Fն!b�����10��5x��OF��ە>}������7z>�s?F����2�~��KpՎo"�n�؍���xe=%�H�~5
��Tg�ѻ����f��PnAg��D��h�iJPku��q���x�`��wV��Y�|��e����۱+;�/ �2ϕ��������?:���!������n3�K[��g���T��CP����(�a����ǟldb�d�CK	�w����kCˊme
�Hg��p���]�����h{({�*w}%J}���=U%X�5�I0�={v���WW��~��K��ɞ�Μ�����TRP0�������sT [�2�T��9���Ш��Xsِ8��
"|K�|�U�X���!D���u�z {�r��o�"�)ے�
�#1��\st��}�J�N�X`Դ�HlS��g�Ǫ�Og�F߰�d�A6�J�kJ����aڄ�/PV�!L�I�V2��M������c �Oǆ͠��k��[R���z��Tm���_(�-��=���X�^R�ne���D��zte6&�����t/C�Pn�|�P{{���N�������'��ߌ9Z�%���:�������p�]gk���c��h_4'���;���-G�;�����'�y��{�:���X������㲩%p�?x�pm	
�u` �)���xz�q���}C֢J|���s�mh���9w������nyzz���o��,g��W1JZ��hEX�.�0��O�o�P	T���4���8+�=�㋑�᧼�&ɽ�,�C�0u�<Y`Y�~P�	�uu}�����5Q�T%R�kw��%ͳ%�}$� QLE[Ϳux����\�%U���): ��!��A|ؤ�(��*eX��W/吝�[����]��ҍ��]������ÉJ$�y�#�D��X6�j����F>��I��
�"j��z���KYv,�gqMLN�yu�ט�Ca������Փ#�jHs�)x�x�uƣ�m<<�~�pԸ�AU�����nih������a���L�pS����b-�(#t+Sר��I������[�x6i���":)�v�n1抌�#�(Q��uS=n���8fS5�����R�"3Y��Ѣ	fBi� ��i����777Gv-pt�>}��Q�Ok]�	LW����Y�����5=[4Ɯ�4����!�ۮ�����'��q��YL�Y��?�D�3�����r� ��dcY�"��aL�X^��9?G6_�>�P}1��F�Ƙ��L��	<f(�z܀�/���M��8J�1
i��k�@6�/�_T[D�p���8�̥�N���������'��ƫ

i�c��QE1�v��q���~�ywP�"�A�+�X��-�/ATo�?�Z��N��>}J��{M5쯅�AIb���kVYY�r"z��_�)���'�K��̚����7�`f
��M��l���\��H-�^��w�Y��g~3�Q�u@�1F@2�v�e��<�!�(�cmZ}���� A����z�p�@ ���ΰ�����%��:v��*j~�F�9>>>���먛���K^^�lC���J�n ��B��n�:��<��/��Su\�eil�3;�F���{��bMK�K18�
S1�C�{��3얠>�]�~��\M>�f���Df�nr��$z���F�[�o�S����OJ�s�&w�q�"jn��Do��ϵo�U��}j##��S���꾍�mц>��3���@]\\�<���V#l玴��\3�E[Z���-n�ט#��D=��8=<��e�Z��\4z�Aqy e���5���߬n�z�՛ٿ��t]Q���Ʒ���;�� �����������L1}�e��H��^t�Ű����� �b���kcҎ�}�&���'xY�,�J_ܴ$�����^�RWܾ�Y�=#���ć�U�Hk(#��r�>!���/�E�2,��u����|�����ɚ��]7h0�."�_)#@=x�v!<l��Nqp��ʊ�[	^qq�%�1��VX$(�1<}j����g�%����lľ�e*?.��i�����p�1K����B�F��!�Lb�?���T�5�f����2�_��E+��� ���:	�%4[r�9��(�n��X3(�YܐY?1#����9*:5;��m{թ��-Y?n,�\����>��P���j��z�@cȵi"C�p>�.�(�����eE��M>Cm}}�F�*yw�}#����T�fol�Y˿�k�t���W��Rቘ�̚n����&���X��d�%�MiI�:�(�]˕�Бn�K�鬾���-��;�B�[K�'�������Ѵ
w4Q瞜UPPn�lO��2�|46	E�Rhi{N)�Q`���IG=�暫�OH��h?ik���c���.T,p��+??꣣#�ՇV5�[�O�^��u��יr��R�ޙV�!}-j s`���t}i��Iϭ�%O%� �Վ�j�YP���e��d�4���p������;kwN�1I�5Y��"j����{��}E�5�(ɷQ���\ԕ�K����<�{ �o[l�9�����o-V��Ln<��噺��>���3��+,G+j�ʠm��yJa�0���>����_:��1�GK.�X�?����j>>�P��g	9x}�i��~�XOD�)w�d�u�s��t+��Ɯ�O�J�����ԥ���8�4/û�t��chb=�mUh��yQ�N��.�s�Ǆ@�rx�%DE�U�C�:?P��:�z���T}�[/=���g06������{��zߠ�t�Q�,�^ZeiÀ@F+�Z�p���OR>�ocZN��'ٶ^nP4tCK��ػ������.>�3~g]�?S�ꗅ/�'�G�`#��_2ߐ���kA����)`������u�ۻYa��U�|i/����@:l9��L�pHN}hkE�cK���ԕL�ϧ^�|T�Х��fN��%M�E�˪1�˵Ͱ��=X<��������{M*$)j�µ�ڢ��
��{�%��`h��CQ�D�P"����� g�\�߄����3>�/������A�Oq`e����d�p�!B\��䩶�I�%B¬޽g�����RG���R֩� B$f=9�z��'��7����k�o�cެsG�
hr��[��_��8�\f"�݀���BMB�E�i����e�}z{{���'W"�LASmM�n�,��8&f��g����/�����s�X�6�*}�A�F�M���� h��o'�{�c��ע#��}��i�sV	�7Z����j��!��A66�|�D�b��f\�T	4��?�8�����%KKK��<������/�P�ge�h�`�/@�`"r��A�a�{�t����nH�-��D�� ]����'�u�:вOɗ2c21����{�o�J����Y�|I,�{E=��Θ�e1\������������3��v�ߛ�� z�\��"��$�����)��(A�+_��9@u��~L�l~CVV�OD���R�v��D0o��[D9SB�'���^bL������X?}!�y!���W�b�k�ɫo�z{�彄��e귿�J�S��1�8n6���ȍh���iK�XT���.*��j��u��%�p�vx�2u�iaG�Z���͉��فu��"4���H�Ct[��ͧ�L+�5!�0 ���֔2��r-��f�lބzj�)?����!���"�&���r5��� ��h�闸�x���:�	$$8' ��]�{<���M��L�e�_��mdyܟ�˛�q\T͵�3��!�3?
�/>���t�����v�����G�=���'��J(Q��]K�yS�^߄�X��x���ߪn�z��ƗB\{�4�������������W�%�����J�(��]<�r����6𡍦UI@����Ug9��~]���9�'����JY�<Pǖe&�XR9��qk[[�L�ț�A��>W
�2<̣	�m��N��ٓIG}��n����^֦�`������&ߴ���A����E^Q��jT�rg�)�l\���58�ܤd��>jW����K�>%Ƀ4���󾆀��.�a��OON�NEސv�Ȳ����T M�T�T8s�Y�5��mO�����e :_$�>i!�,&��h�:�§�xCY��̘N��k�J��� �G��q�0.���>LC#�T߀�Or��5�.2���ԃ�mx���]i ��N�)�.7�ME��T�m@��S{I*��G�h���MODYb�٥^�����k����Alɪ�Z�ΠRP�D)�?.�g�#�|�sGߵ�`&�I���}�{O1u%gE�ˤ�nYW(�~V&m��cnR2y����;�,�9���ϟ�A��Hv�;�Կ�mz�������Y���?� k���ǑO���n{#)Y��<���l����j�7���#�üV�U���~_L��Ҋb��'Y�����7�b"8��H��q��Hy�Vg�����mm/�����O�ϛ�W�u�K�r�����%p���;V�x�bM�]k�vj��+��v�����0KNcv�����-��{�!�趩��؁��$���̆k����coį�ZKب�� �w:�����ְ��x�����#��P&��\����K�f�������M�_T}D;���A���.]�̾JV�������F�YKM7�-���Ht�E�bw�wa�uO7���nE�!	U��1C{?�(����p����18\���I ������\C���~���X��߾���@b���^;X���Ő�f�R0��ncJV,��֘?B�����jhj�$��Z��]r�Y�篁&4KH���q	�������� n|��?�~�Tx������'���Gky�e��u��L-�q�3!`�D���� ��P(T��9��A#��f~��R��L��QqzA&���� a��=�h�)Ei����$a�R�5���'���o�~�����ǖ�8χ�/�׻�P�7��oW^M�L�K �b���OѳP������7����F]!��=�~:��8�2㛁N�� �WR��ߔ�*�J|�Q?��8�GOњ�W�o��N]"�/�0��g�?�Q���S|zݳa��mw�|��c���?:3�wJ���z�0��\~I�w����3��,��a�%�����M�:oH�B\w��W^f�,c��t��B�%��1��fB�(�/�X@_�JA��8�]��C���m�����U�М����<H��8$������^�vI:TD���>�������Q�L�)c�-Q����$A�T5Y<���� ��J��QL�j+�`l�y¼��@l��t��=5I��O�7G�y�Q1��
�~��
i���B}�����)�-�ӯS���*YX���xC`L&���J�oBΉ4�g�$jҥ�,�[o��R��`]�ߔ�e	��9����m�����}>�?��?QjXR(��m_�|j�F����#\���� �"�$	:e�$���W�S9b���ߢ��.�����D��3�M�6E�i�C�/�E��h�tC��Dǘ��I��Gb���c�I=M��<�eX*_%#]�u���l��P]n����x�j�TL��[j�kG�]}�%���W�1?.�,����W��:`�G�����������IU
���E��������������dѷ�y������ӭ�VT2���-��a��1�(0���́P�(��ľ�R�]I�!�=��x�U*�ao�TEw�?Q��D��*]	���G���t
���*�zv�Ft�g�c���ʲ��������C��ٯ��#mÞ�:�e�bꜵͷ����(��H�#]£����h���8D�'m�ߵ�u�Áp	���]��?m�r�t]�����q�y�o�w�v̼�D�R��_xЧ �pZ�W0�x�Y�X��KqKL��@?�:�9�|u\}2�p��|B��W����f��A}_�c�|`&��Ȳc�*��s�#Qm~/厮$�}�i�hN}�z=5����r�R	D��k�����.d�K��љ�(���A��C�-��k����U׼�-�7�䪂��Ԉ>��Nc-�>L�Or��yty%J���/����$�⨩�ۭ��ж;��F�,��	yg����I;zHGE�!�6��L$�[^�l���MܰS�y��Ĝ�t����ջ,���|�=���YH�44y�)i4ߘR����H�k�7����fN���'�����8�~�I�|�%�Z7��bʥx�4￟��TD���E!4����{@K�q�]��`�.�=f?I��������,:��6���E�=#�_�oi�<�yM+߀݁���N>�xZ�R�6�~Z߇�"�&��?U�$�+�e3��
�,9�~��ZmF�8z)�6�c��7�~y	9V�����#ԃW �2�Kj��9Й���z����� :t�)��~�Y��t�]���䓣w/�%��0��:��d�좗w��q�{��J�x��1--]F�p�����&p@_;��b��؅�Ԡ���;7x�����>��']�!
�������yܮG� �^���*��+U�N���y���1����eƿo�5=��� �@0Ù�4ٝG�4�M��{���O7|u�������y��e��<�[��-��5>�MTEH����o��tj;��)���ǈ<�x���/w�����9���$�Ή��%���?$�>�F�W3���{��Y�?\F��g,�p"�+�JP�v/��J�]���+h%�f�~�M9mi�B��
�{ �Dk{?6z��咈i�5p�s���r_x��F<硍���b�ז��}��'������j�@����N�nDJ�A:�$��.)iP鎡K��n�.�~Ϲw���y{-�b����/��C�g�~��!�����]��ihr��nqa�*r�r�-ɨX^��-��QA���ֻl�ண�`>0N}"(����t�#G�f�������w�c��,7�l@�欲K�����F	���NN��%�W&���w�v��F�(����B�$�h�}zPC�73tu�A��#�U� �}�jJJ������)R�&�i���O � ��Mؠ���_0P��;���fH����#9.�ȈEg�~d�����|���f�c�2G��a!�
������������v:����n{����$I#_p��S�=&���3�I�������I$`��wO��cN��e߰�z�C���-��*zX�J�]�KаJ��H��6�jCt�ށ�ࡋ��B���y����"�Ӕe�n+V�H���+��wॗ]X�W:���Ij��u���7���(�Gi S�D{cIٴ���
��<�ۓg���|��V��%�#i�=�[xt�}򶀜iM�ۊN�;,�#k��ԭ�۵x[z<n}��`~٣f-��i���^�Uk��n�M�����&a�B�3���V�����f����*�ǯ�yϻf1��1l�۬�4C��g�[��t>��*R�7�t�$/RK�[w�1���1����x��Z�Ⴆss�b�(g��6�v���B�W.Q����i�8>���3d?pr���Y�xR�_�t�@#x���J�5�ڬ�u�t�����衟pڈj��=jd?�0�]k��'��LjdE�NYn���'�6��	�M]��˯����-c��e�����w������6����ma[[>���Yܟ��$�ʾD0w�SɁ�o�o����}��Q�+�v<�^9���`k��[��5�.�i֩qڛ��
A��{C�A���S� q.�kV���?@ ������U�C�=��7���U=��a�=�Oֳߊ��YL�L���vr�B=�]6kϡ$�u��ZX$�\^�L�-�Xԧ�jC����# ԩ��q����#7i�|R��'�3�qZ��!�F���,�������Z���Չ3�|�u���ڪ�o��N~��1����H��x�{���T/6���o�w�O��l���GOa������3���_ ж�%�5���
��Wdu���j�� �5����j;���t��p�se��N(�?zz�K
A��l�#.�1���G�V���^�5��o�9�s=x���wNo-���XJ0����@C_a]6,��O
S���ΐ�k\6����K*��w����5胵�K��畷�f�ؤ���^�}=���?�ަ+�mu���~� �9�`+�;b�m��<Xk+l�({ѳn��`W��ԫ����u�X�tHa���-[�@t�mrZC`���C�x&�S���k'IQ�/�\_(Ry��7���n�d�.ف�y��kC��nļ��'��17!���#�T� �X�` a�ήx����VCk�	<ͩN�]�����*G>p!A���
����@IӴ��f9i��Sv_��f����&�KY��תAϹ�q�׃�G�?�Z�:LaM�aS$�\�&9�Y|������-��_��o����Z-ק���QQ�k9v�cw����~}���G�]�.���q�K)E���j�d6�'s[��d�ꋁ��l�������Uzi���Ŏ&�@����b<b~���6��5z��|�5L�e\�a����s�'��o���Mͷt#��;��eΐ�q��� OmN��;e`�Ւ����ր.�~<̏P���7Mܩ�iF$�vچ�ą�yC��v�!�(ۨ
|�8��h�����~S�`����t!6u��Z�r
f�l���0�>��3]!�#R.�.�g1i�˪�fr�$L�5F�,،%��,��\7@�$�ՠ��Ӯ�)��5ev:9	�:|R��0Ĭ�V�L%o��ĆsI�C�6���z98g���
IA^��R�z6��y/6q��Y+P����1��.�5/Ch�$��EJꛤtY�su�m�zGj��ѯ�%��E�Gmq%�uL�w������nK�Mx�r��"Dj�X�K�|����l�:�12���a���.j�@O�Ɵ�/�h�lW��N�uA9DӚ7�˟���Z�K?V�aI�M`ध牛����[�P��<���y5.-#1`䃲��Z��AH�A�'�����05`Q(IIeͪ�7QH��L��.'���!�+J�{���-�/3�<>K�I��QWT�r��;_h� U���Z�����6�;uB{!��h����\Iۋ�Qv�E���6�g���AC��2F{�@���$�'�̒��+7�IB�@-�_&:u�}����#��8�&��Q��k|\���@@r�d�G�MA�rT�i�Ȑ	�oQk�=7J�����tV��}bu��r��J�������/|�Fn�#
-G�������m�e�w5s�H"D$Q!&�f���*�F_����u !p��?*���vu =�y�������w���3�@|�)�ػE�x��	����d�n3����R���޾u�gdP���(Z���<u����5-�v�K�i���g�|) �C:.��gD�d�l���S;]P'��9�'7#V�Sw���#E̓���,�)E�@�����6,V7y�����-Kܪol����j�Bk���q�r�ڃ��n$�P�|��i=]�w�-�;Y�u�g��х�o�H$�yV���S}k��o�9��|�n�,9�� �z��H
�m�}W�5wR�	�U2C�Ѻ}���,�#p�����M��^_�٘zV�C���tժ���6l!���i�شa��R�3
��!D��������p�2ٱ`��c�B�"�,��}6|=�9�%�Π��Î�Bcc�A�#�)���Be9�?�Vm�&��Vb����%����k����c8���"�/?�gX��
�V����Ù}�:�� ��e �p*���c�ܞ��vA���i�v"�����K�</����[ή�>C���Z�����;dG��k2����ˁ���=9�-l\~~D79Ka�6�.�`\�%�W��a�h��
�_Ԫ�\��6�=$�#�G�K~3��\�ռ�V'��C��y�!���-����H��60X�� $c -�E��r�FE�Y�UVкNtKtH��Y�Լ��Zq};�1kY�!��f�*xa��AB�C16��y�?��}�opJ�������E�tHWw-Ѳ�U|&-��cm> ��t��[�h���F��])h��N�^�b3�˲�F8��ϐf��L���h.�]d���g4�@�
u��4�����+���J�r���^7[��Qtm��&�?H��Έ
�Q�g�O�J�c9r^M�hK������zK��>���n8u��59i����Q1�4*-�>��K�*L.�S��8(S�4Ζl��B����1�C
�;"̀屠w��?׃���B���\+Mtu�rfs�`��l	F��F3]�x~c	�͟���.Ε���u��ze�CEҺq]N]H�����������n:y �a?k���b.�.����q(�!	���8��^*77�1:h��r�)v�[QQh�6�ߠn�E4~��t��! ��+=��竿�GDlj��P�}51-�&�z76�����G���%)0��nbo�qf�����[)_&8S���ȵ̳�*�_��_�%�	r��$�֞5��|�&��gHwH�,8ޝ��	�U=�*�}'Du�>+�E"��
�b��˾��"X,ov���	��e�>o,^{���dB93��SeQ����
����Qs[Nk����rH�'OO�I�K���({��Rƣ�ImU������_?�a���,Sٝ�����2�Ŋj���O���!,�2�������Y�����2���f�a�}�� Е�nU��o�3`?�7V�.��(8�c��n|n�R���ᔕRG>6�"̛�����IC"���>�JJH
���-�Y�ƺj�yc��3~�fE)������];���K�*�^He��yV�F�u?0��?��na���v`t�J�k�g�"�.��lO.��A��U����;�Y��O(c�ȯ��Ϻf?kW�Ę�[�s�ur�F�[EG��8��Gr�"q-%8RIr�W����+�W��:SA5�B><
��X	k�X-G�2|�`=�݂��(�Q�$N>�ѷ�yִ��ʪ(�^����N���HZ����qq���*oo��Hew���~�K[3��Z��3�Aↇ��Igb��~�vn",����? J�A���Ȭ�L&��"A ��l\?���-^G��w駨��9
]� ��C����:��
��U�7�O�s�F����, �luW%"��]b��g��Mp��W�u?�δ�\r�0����I��hJ���?�����A$-hN����cJ�;O����PT�����/�m�6]މ5�9gRLJ��K�gi#]ZC33�/c�B�B\Qd��qf��M�� V��z]�EV��
�F��u���)6��נ��}3�r*z�C���V��O�@2�Z:�E���v����A	'S*��?1׈Ӗ�ryj@�SL|��bE[�5���12��}�aW�+�$�P��hz}�~�����I?�����O�������W'�n���|A%�$֓�U��D�K�F@�*�X�u�(^�R��TH(S�˹�]���M�G����(n�E���}+,�������c��ɹQ��ldč������\l��q�6qwR�v����Je9�H��h�k�0_���<F��\�o�-�Ln,ԂF<�r��ն��#����*��h�n�!�R��C�����]P�
ذ�&i���ۂ4C�?�m���S��*B#Տ�"ʀ��3���)���8�S�W����}FmVhHmT+J�l�@o�lyJ
��k6�����F="���q����v���'���c���N|�����k�"�Y� �OK_9�A��ϑ@�n�D��@�-^� �≀�����醽�w-��_`DL�5��W!_p)�����mH��
����/�\b�Q�+:7 4�y�� [�7h�}�;i�>��Skh�2 a��"M�i�5�c\"©�%�*��7�lr.0�rX��g��윫M�`y��<9A|s�=@�f���$o�&��JbTi���[Uh����Eݢ$^�u~�"��ԲS��6n���w�ov�=�RT��Y� ���Kř���St J%�:)ޑ���_d�jd��W7x������:�ʤ�(/�-�q�&ˬ�LT=^JO�Z7(ӆj�)���<�a@�Eb��E�����.�=?]�I�׃�j�8������[�䔧{�檀�~)��B����	�%���8��=�Q��:��^���O5!3Z������=^n�p�E�4�0�& �.���_�Am$����3���s����������Cqj��/A*���3DNb+�w1c� Ӑ����kb����Ds�H�,�;4�Y��[^l�M%U�`�����MA�ԝ� f�<3��ӣX�b+!p{E��� ���~��,��Y.�I�,�?�w�
��>��.�8b]��"�ӇψF�*���s���a��*��.���fԩoW���U�R���*��b��VԵ�a�����Bi[^'W�V#���oe��?����ݲS�R��{�8�P ������(���3h7�F��+Z$��P�{�P3��gĚ%V�	��u~@�����s�X�ĸ/C����a�!^�UV��F�$�eA��<��&˖S���j�����AbB���2���h�	�Q�YFQ~+����,�]9)����NV좆U�7��� н�R�V��||�!�U��ݪ� ��O��jG%f�i��25*�Q{�k$�8S���J^�.�u��9<�aJF�-�L�fX ����Ã��LO���sܢ��pUM��ig�d0~,�@\;��pC���u��%S��^jclSM�!N��;�ƙsF΁�1��o��D�7�`c������`���{�� ����M��Dz�O�q��c��CH7۟Yo�ΦC_�#�p��/.X�x9�� u�2:�Z�ˁظ;���L^.R�7^������n�����e��F�!���.0�yE΂�c�����
�O�%�%��7�E6�אzxr���k�(P�y
GA^�RRFt���;��`2T�{>���9{ЕF��g��%����yZq(ns�,�+���T�=
$=@Ϡ��!j?��5ө�$���CRT�3"^3a?��rY�e,S#/l7�"���j+�Y��Y�2��-��ma�7w�>�6Q:�\���c?Ec��( d��TT�L�Arr�z�^S�(Jؕj{E�\"�!kjf�����X&:Օ���>!Ln5�J� #'�j{�P9�Q�Ms��l���v7��E���E&��	�ׯ�G�:��>3�)�N�[�yCy�Lh����.�`����z�@%�����"��bU�dgS�ܟ��B�b�����;� �.��������	B�+�W��fTä�JO����: � 7��~�����x	m�u�ѓ�aou�����N J�m�ی�i}a��SJ��nϬ5�hd��X�|��YG��T�]\��vX�9�tv�(��9X@��O11w|��h ,*k��8e\��"2I�S�a`:�I�sSO1NԲ��T�m�N���Q��A54\S�[*Ns��.����������e;��͞vn�"z)�_�C����a��^?�7���X��%�
��m^��vR�Y��h:�"��1*�YW?���帽�z�̪I
�~j��D+��$�L�2���Luk��g<��lӞn�a�O�#��O8�F�ရ.`�o���+l��� p����D�1/�M�����1���g[DGϨ�Ef �8F�8W^b:|a��l�eғ�@T��� k��-M�.�����_��G�b��A?�|�-��Hb=��;�9�;b�IQ�8�!�j��
�M\"h���<v��o݌i��$�p�^�I�vcS��n��߲��F�&�?�o�&�ʛ�4iR����9$�>�dUVeg����@��V���?Y����d�SL�*�XB
�7D��f�:	M�Oq��BTON�˔�<ƞ�Ҩi��4�/�|-'4��)�)6q��V\~5��9��M���&i�����Y�VS�(<R��!�u�����i�*��ۘ�u�͛��h`[�~���F#�8�4P��e���I�P�/F:�T�냷��!���.-�`�!�g+E�-�Aߥ;��#g�ò�;82�=�$ę?�Q>ڒN_��I_]d[����!�2��F�y���}1�Qb�����M@�3�ګ���m��uy�� ����O��
!�u~v�����t.Y`�_|"=�knG��<m�Oe?����OY���$o&��{�iAǜ�j����X2���X(QmiM�FeZ�^�͍���Lb�U3X�gWf���M���T����CI��h�f��T:)���V�7�FV�C��ariN�.�p #���-倝�}M������c:�5n.�[|Ӏ 	�HhՁ(��DZ�9V3�� F��"��s�*u)L�>��G���IЅ�l"e]i5LR����I8��Z��[q�ht���/���>��b���[�^�&�wv��V��pK�a�}���������H���� j�DT;��Dv�\.��#*��6�����O3�J���.zM�T@�LW<���=T�rr�Y_�k����r�%(���f';A�9 MQDØ��bV=9�4]��y��M���%������ �����:�h��C�)gَ����"�߾}���5��BP�~[�Dꪲ!��n3�R�f��m��n8�k�A��E�m��T��0c��Y.���0����q�$p,R�}�p�z$RٝTY�t���uT�&�+G�FA=��)����C<Q�׺)L�!eP�JR�ь�s�^��n�"= %B�r]wd��t��C�u�xL�,:R VU�u��(�v�H���yX�w���8�9�'O�,�=ߘ7|�w��,&1�o�IX��N�ª��VY��?RS��|�':�Tv�n����󝠍�`�J9���庚a��H���pPv�w^��vj�b���	�}�s��Y�=_i��D.!̨Z.�pɟ�ǺdVTz��z{��*			�GmQ퀉���$�OE`����w��Z����m�*��5xP�H�qW���!%!��b�ҬD��QQ���y����g��.%�ѫ�1:��e�04\���w��١�K'���+I{�\�+�@��EV��ә�t:��;�d^�Lx���f�&�½�BjsGv��1<+�zJ�(�H:��Cΰ���$��n�kzХ*T�@�F�v^�מ�_K����e�u-:����Ϸg/xU��/�Ӭ����0�
f�ڶQQ:UJ:UW��5�N�	�"���o�R���U@/m���aOô�5�^zk$�bd��pƹ��h���mY���{�L�J�,[|Ka�MN�2� �[��P-J)�J�©�c�\Y���,���:=��M2�J��@���aE�	)P"�(~b��ō�>��N��#8Ra��v-P��95�֔\�5�pɫz4������u�)%�L6��`�΀$�ǋU�I�x:Y�� Io���-Ʈ<F��o�H�E󱭹�8~iY�"�.)�@e,��p�ݘ8�,��L���<�E2#������f��*g���zb'F�O(���ʴ-��]�G63d����k"C��\�瀰w���z���+\�:��M�(b�d��ac�;:���K�^���^�آ�t�,'�-q�Ǉs�UqJ�����1 �K�rQ����-������P�w
�]�q	���^.���@T^nq�-���Ẃ-���r"!"!����S����xW�2�_����HK��8l�Nj8'�"*e�O��YT����S�
��Ҽς�t�%��ͭ(�v�"�N��T�L�� �4B�a�k�@֩,P���`EiB.��e=�;�G�/�'m�𕨓�EcVQ;2�7��a��kqq��vX!O1��D;��lc�Q^imĩ�q~��U,�}w��8y���s'T�4����m�`ۢE�C�E�o��U�1��KH�m_*�����ל���̛�^�j ���������W�wuopODل+��`�R�"��������6\--u���M���?V��@U���&���|*�]�a�LR��;�����+��5HT1+��i�U��"]C+�8f/(�!��۷�V����a�|��o�Y�u�b3IL$�����S��|��A�K�yM�^�˂E��
���\�W�ϼ�sd�W�:�7��5h[����e+��=1K%?/��n����������y�u@��E"��̪HAQ����x[o���b{��J��;�v̴#��
ڬ^7���2�α�ޜt��.����Ӧ6�<�K&ʀ�;'�v���7�)��9�m/�Dt��D��g��=ݢ��J�c�%p��w�����+,� <'�2c�n��ca�ÌR�R4�rU��y,Zh���6id%
�(�ػ�Y� ed���飁�A$�U�=���#ˑ�>���U,�s@�r�l��c�N?zn�4z����o�KH8�<��H�qϪ'���"9�قR��dF�kH3�G��ɍ>\e�m�>C=�q[���E�cu���z�'���mF�uD]FǠѲ�TU�@:�����s��V ����o	p	k�������Ή_O�fM���y�H���Iy	� �N-�.���P���%&&��&����X4F���Q3���5�w�/E��9�����N���;�;:�48�F�(U���_c���$/E�G��j� �oM��Fx3i�
����=ޅ�7�����DHW�Һ����,C5k��v�wA�͏P/	|���;�j�}�!�k%�Q�[˳%�������A���'�T�
؝W#��{Y�?���?����N������^�F��۾����4c��|�l"��%k�橝��~Q'wa��1����������]��(ˈ;Z�� a� ��V�_7��r��z���!X(��p��8B7�¾��w�m���9��?�"��:d���赑�)�����x��I�����֞5�����Q�n����>ť������jֵ3/JA�d�[� #1h�(��~z��Խh2�R�ĞZ�L8�	=��&J�����%�dw�	4 �LF+�p�3_�|3��"�a?XVb�Wt�����S!]�SD`�M��$�]�S6���qF�(�7fA>$/�#�/'>�Q�y�I��3�7I�"Ў���P1�Š�u�m%k�2�� �����?i�Łُ�Z�N6�����4}0����"Y��B~Y�:��IO���X�|�u5û��<h��X���х��j��+�̪;�o��Hq�^�kVװ:���5���e��,����9bco� 55�doxH��r�DҢ f�9��!	�����&p�<��D$"���i�(�?���KB׌k짐���[9I��2��*��Jk����5꽄���-��F�G�y�l��v=!��Yɡ�_�_���peNl���\��0����юd��A���]�b�@����C�+�d���bQmu�9�{��s����X8I9�v�5J�;�kM��3�V���N7��m�`xTά�ss;�m��D�����S�X'���������VԣU�]��U���D��1O�e��l�.t�x����2-�79�����5[ƹ�L���E�/�pU�\[���#Bϡkb[9��.�����F�ͬnjƚ�qѷ��K���hn��%(P{ �r EY�
�����$Zʬ��»���'�}�k^(Hۯ}��gH�V6=�]9x�]ahL��Ǒ"�}�5�*�w#��s.�|r�2##�V|��;��D;�~Q%5�?���9iXB�(�Ū���3�u��)�v0>����b���C���p�V(��
k|�[V���������K�Ynn/_����)�����<e�Q���	34�<f$�J���	���bK�g&߇M�kN`y�i�pL���I�j��{X߄tF��¿��U^�Đ/��;�����_*�]z�q,�ߒ���4�վO�ir�\1UC�(:��P��x��tRqV������[���Y6���� ���b~���f<�!������Su=����A۶�5��㳵/��{�'�4�S�i=��M*��ޙ��٨�>�������b�
a�h9x��hf�C2��3�=�%�
H��m�:E=��Zr�]�_V����󅧫VעPo-}p�fg�]YANeEP'$���$R�r����p�t��=ȑ��oM1��.V�p~DIU *X����p�v�{���mE+��d9�'��:X 2�ʩR]�C�+Ę��j���7[S������[�����]������*��d-`u��}wA�~�N�iF��x�z��Υ?K�:�`�<�f�l�{��(�NR���Rp�,[�Ȗ�`8��ߵ�MFVy(�7Z����(���j�N���w��7���$�hy���`�e��W�l9^+J�wTO��d���F=1�0�.��R()�Oq ���i�I�P���Ѝr��j3�1ֆ8���B|d4X���{�٪ �z~�l�#�Y~~WΟ4���/#���YX���T96��1��	~�n|X�)Y�q�2qއ�0:����IT�7�I�O�­���סּ��>��،�3������� �}�G��W<1\�0�m(��1լ�k8��}de�2$��y���g$pݙ9�� t�8�8,�;���t_W���M�qz�b�j콡'y�1�Ą��fGd�_��8�Yx愅@���H|��1��L�4\�`8���)�����}ڲN�wJ]k-�?,�e����(��:�?hڤgp]B#$Uҁ@~!��Ɋ��vL�o�W4$��Qh�R��r�n��hZ�+D,�C1�ȉȿ9�{�����<:���-�v��
NJ�Z�����B`������a�"����?N�1�Ճ���=z�kQ�ʯe:����6�:����/���'m$j�F"���-�ݺ��!V�^Z�LU��F��i�u'�8<�%���ɷ�#HJ��E�ܔa=9_��0VII؛y����
����W���s��љ�sz��L�q��ć�����ry��Gs?�%����.J�L�����`��݄��Ʃk�D�e�R�:=ъ�z���ҧ�f#^~��T�4^��{;������Ԥ�����YjUč(�����y�?��=a�q��,�
H�e��90�v���d�~ZKx��4���? �y�c�r�\�󓓐�l�$���H�*Ec����R��4E�]@4�?l�j��x}{��H�[S�$�{\mra���s���P�x�S���z(·�MHe�dԢ������)�b�|�,����A���Λ�aWX<�Ly5?.x�<x�[
5�cv�9��G�yQ��hz���bl8�P���������8�����V�x�tB4@����D��{�(����} ��F����ɏ<K��[E/�0)`m����߲MblS$x\d�Kd�*H�=����L�pZ{=F_��C�o}���i�]�k`�)�F���Lś���ϐ��:�tׂV2�7v�N�$o^�l	G��kм�������*���D���gΚ_��.�;��܌c̼���t���tz|�m�˴@�1��wh+�=�}H��v�i�X}�=YN�t|w��5<hμf��&��F�qz}��ᾛ��!o��lp��kUK���W�^�L~�T�:$�*�m.���h���*�\�Oi'����: ���&zI�+u�uo�y�z�]��*ް��F��n
9��j������� ���|�	W8j�T�Y�D��:��lx�Y����Z�K�7y�d�.o`/��騆l�N�}���|�vT�o�m �)�T1wM2�dhD~u�ov��R�����{��������Q�n�om��\�e�/���a����v@*������DBY��Ҋ�|E�dC�� ����z{/�~6a��sF8c�d�l�\�Q'�ZBt�>ۘl�'�$���&�ۻ�mq���ٕ�����u���7\���Ѱ��?�����L�V��2�g�M|������Gb��bB8�G�D���[J�@��Ƶ|���z��BcDcJ�o����Ki���ȡ���������\K��CD�\���f'���kz��JM������P �2�E���uK�����4Tn4�ς�Ӄ��&�^�g+�������*������� ��Ij�������G���a�&?PV���llh�I��d��@������%̑eqa"j������R�,�	r��|�qN�����B��#�1t�M�n���L�P����q���t݉��}����t � *a�w,a 1�Gs��b�|`��\�T��ހ7�n�CsMx���gz�rV�1r04�i��_�+����� ����J�2� �c�n�r@�y��-�`�;�0 �C�p��hS����W^G���4<��Ԝ���Ž���Oe��F��G�k�֒�Q	gN������g��qvʜm�6�!`���1� �,�&�X���-ޜ�^n�RV�x�l����%5�=��B?���֚�8�_Q�@=k�����s���$�g��	������[gw9[w�+��g�b��F-��<�,{Z�>�������X3��\��'�\�:��ۉ�0"B�?�EfN6T�؇;���^`���?�^
��̹��H[��yB�E��j�}ۢE�5��,eU��H@��ms��uE�7�x,�0������-I�h�[͏�z��a������zBQF	�Z�!%%�k��Y[�!�LM�l�~����������P���A������U8w��?���Zmfw��?,}9���(�*�`�Pé<X� �[�g^��wh��6=e�t����I�xi�2�S_ĲQR@{ a3؜w��+�-&"7��&rޗ�Hl����*aS�#��1���cv+�� 1e�
�E~�����0魧�a���TOf��*��7�ɮ:+ޒL�����3o��r4M `D��)�������j6�,��-�Yq/�[�*өy������AE����+!�����}N�&*�A��!�����]|\����9\�I��s�
�6��Wo����t�:�~u�e�-�:��8��;ě��<�u���q�]x����\��y�T߹���s~��>͝�?9�J�er���&ˢ�,��I�3��ܲ���p�������'�U\�;�f5^���&,e��%�iO���",O%z�?����G��j�ʘ*>�$���̚�oyC^��d)�吥�����/my�����q�P���a'�#����ʼ"��Cs�hd̹M�v��YL�߃����%�'��pҷ���n���҂,,T�d��Ot��&�&3G��k�f�i�-��q���`�k�ц��Z�ѤD��+��`r _����\d%1O0���Ja���,��	���w���L��ة����Z�n��W]�5�RAz�d�@�e����e#��s	�J�8�9�gO1Q��"��N��[}��fu����ص\�!mѳ��բusq��:VD��_��ӏl�������_����-M{�9�_�o��Vɤ�)J�5���M���:Ϗm=HP8m�񣹁�pb���C�CI!���]��p�t��z>Q,&���� u�|�m�Į;gs�a廬Vr9kV(9K��WX9��1CY�7��7z�5y���������-�����c3_�^!傢��l)\ՏH���o蚅X,XH���W���
��^|��m���8%^p��Lbb����wl	�0�U�FO�y���Q^�����'~u!(���o��G�[��s�e�+9^�/C��c����L�E�f�sS���e4��GF@J�(�1-���Nw��i�]ԩx@��@����HT�g���O�N�g &C����3dK��u�����8���&����q0�ǰ�Ecp�F!)��=r��u�Ҋ�Ƽ������0 ���7#�:�+B	��/o�,���W='���^ԟK�pTf�N8�Wզ�%6n�!�te�y��r�rU �=�'+��B���G�D�)a�k�e��X�r@-���|̲��m�kCU��ӕ%-Au�x���칢f�
�F[ �����1;����_���ܖ�����~yZy�#ֵMc�A��e�'������)�~��+��t��l����'	v������0f�]�x�K�x`�D��r��j9��� �:h�D�}��1TU��e�{B$��e��1�Iy��O�J��+�#+%�'��v���sc5����د���=��B^��K��C1Q��=1��B#���ar�mw�d��K�9��=)�%R�+5�ȇ�dv�D�\��Ӎ�wG��u��<���!�7&����I�\���bz��߅�X�C:�X������q���fK.��;�s����(}>�̟5��~��z&QHns�P�:�GK	�D���]]49����E/�R�H��o;K���gS5/�z�
W�҄f����kO5����"��C��C�wT�Y�u>M�+�q��v�ϫ�G}����	bR;�2����(����bP�t<w.�=�n�?�hQs�9=�||��sN�vp��m	�@N�j��tDD,}T��n�`�C1����b���z�wb�M��^fL+��������k�L j��u��_�*���b�3���Sb��]�@���u�Sm>B���'lNuX���_��b�?� �� �N!��	��ڬ�X���F-K�`Q�:��D*�U>���z�����h{�+F�Tr�憞�v���=��p%����V���Y�'�$����͆+�Mr��h��[��$`V�4+�V]��������w~�V/ Η�n�*-�o���[ͤJ��#ay�����9�.�#��e\�pf�8�'"ċ�-�+Ec��e���ܭ#���u�Gal��e�Z�D���ҘURs��8��+N��k`ސ�\!8ն��F*�>d�Y�\;�ȹΟ�)�{���'�.�{|��m�j?��|xXQ>��į$��
����`%ՒOӄ��*㞺#W���w���ކ�@u$珌��T�ޔN�����H���_>q̓����9^�'�cOL2�����-ɯӡɳ��'NP~��`�c�l0ANdq����E�����K*�t3����#5��m[nޗ����n�N���9�(rZ�(�P��O;�Y�C�-Gj�=U�����O��;��uq���XJs�a�^�Bu���0uTO�iÇ���{:-Ք�r�})��ݠܳ��֧����h����SW�I�6i�|���k�7�*��w�\=���@���߰���8�t�罹o��H��쯗:�{No/����n�ot��1X;� �pQ�;� +�S;{!��s��@H��zy�b���{W'�P��f\q��Los�^�q�DB���ch�Õ�w$v�c��������T�-3��b���C#ƪī�y�%Q]�d�̹��+��*�̏?r�r0t���n72�M���zG��<�z�ُ���k��)�u�Y��:��П�t�כD$�%"'"'��]�K��faa�~��(OU�t��{�_ټ/6E,!z:��*)�4j�ګ���%��f�J��i짪���2!�X�g�Bg��!��T���%Ҥ����H�& M�*�}U��^��t�TJ�Ho)��Kb$@ �'����������X+�s��3�g�yfv����'--?��mB����2p����������Ͷ^��ٺ��K��n����������VS�s�7�v��zwW���M?��8���q�fx�����������iy����+!9W�b�9�{f�����0>�����.ɘ ��@D�"4��/��*ReD03��_��� l`��������l/g��8�x.�k ټk$o�y���kbz��p��)�������v�+?O��O�+o�$�e��Ӆ��T�N(5�W�'Q�K}��'�Fs�]T��h�����q���ԝȻ�R-f�M��N�5��>?��X$�����B� ЄXx��$�2�v���vǜ����	�Tp�0 ���Ѻ{r�x2��&iȊ;�tFҾҚy�����s�����o�υ�ভ+<�:��F�=g�C��*Yq�%(���}�
z����&:vu�HGvH_�iI�~�ѣ�{C� �w����Wÿ��.�����(�e�P��'˩�C�w�(��쿃���;�J���Kw�Ԏ��3���e��z��ǽ@@���Ǎ
�;��rGOO�Pz�"��ܧ�Y�:vf�����'"��c5]�����Ӷꈊ�$�,�oQ#4���O���a���y�wM_�Ѩ$��|��OD.�l��ꢑ8�ɰM�.M7��5V��N��}iN����lL}�}��`�o�T�^G��ฺ�M����p�	���y����zF��TೇX�j��rz��L�+Ǣ�K�/�1�����X��MU���/F�`^0Q�\~!�9�κ�f:O���F'6����.��� ����R��sz_�E��� <��֭�l��K�PJ�l��>����1)x����'�\ Њ,���@kDV��xo��%/[fLj��ϭG)2��r���ǲQ�F5[ӛ�P�x�a��'[�\���x�w{��B�V��(��ٺ!q�`PRN���>я�n�d��O��+f�`�҇�WJ<�Ҭ�ܩ�������YM�wë*��{p?-�ܡ׭�"]�9ʚso������&�Ӥ��l�Rry��rj,=�Osi�+���e��<��-����٢�B�A�Tt���b(4>��ڻk�"]};�����{��������Gn�z<�d|ʚ�<t��$�[��]s�kj���2��a�j@�i���Q|K�]�H`iǓg��Q6���7����҆����<{�	o�'��a)�&���V"x��xH NS7������(8�c���Tc���Ʀ1@�㠟��*�cW[hs)��`޹H�s�:3:�?����o�+I�u��<���^4�&�u���=� B�L/ڭ�0���Km򱡛q`�}��:��̒�̬�kh�r�7��֏��vB�����wi-\�F^���c�X)���L%��ߩ^s⊺T��O�[^o�ζ}��[7���E��9'�q�M�c�Gl,���Y�U��U�)||6�#m]1Sͥ�v���|�?���YXJ�U�r30\�����֝6��q/�_.��h����÷�yQ�{��ĩa���C�u�D��B��A/�����f5K�*�ڤh�W�HqW�?�r��	G0g<��}�a��>�9;���V�2�_�;�x�0�,�I����F=�]9��8�+�$�����1M�t��*�E9<Z��ĕe.t뗲Ϲ[��jڪ�������������O-_0Y��J��c�@�;,������K&��#�P�ke||�?eI�C�+�v������u�'wZa? A���_�d����I^Cq8��Ԩ�}��\Ɠ���7i�s���?���\�O��̞p3�3��ٗ�����v��@�d.��ewNdV�lA��`a��N_B����9�m�ko4.pr�&��ݒ�O�:�P��iŗl̬춚���5��S�`�����Q$B�X�zO������/�[�w��I-�lŉM�c�~Q��L��`k�O�m�w�K��[�̵9��.}�*Л�B<��	Ú����x?~q��/^ʳ�	����u��sd�ffڗ��- �d�����7Q�i9�qDq��z��Ğ ����/�?i�M�E~��^Z>_���/�/�3���SjÓ�T�����Hy#��d�3Uں�俷���R��}Lw��`�2HŽ?�0�|=N��[8�Z���.L��A�#n>ۤkB�\?��$]�(�g�#"�[�F�6O\���Y+�b���,h�G_�
T|j7��;S�?�4���Yw�K)VZ�n"$W�?u��m_�&..W�r�������G�_ �*�ڇ(C�,���;x��b(��!L�����џ|�n��V�U���Y6W��ۮ���Q�L�}��!�-k?���jHf3o$�Ejx+p;矑�������3��$N��������r��G����Fo�G�%��40�i�cӥ!��J=9t� ����-�t�c���g�I�n|uxvu߫�A�-�+�y)��!�Q�V����-c�S%e󁱁���Rp�ز�ߏ��S�a���YB�f.H:��U.ع)ӛ�>2K��LC���f��q�x�ލ�_h���A�4Ҿ��b�ld�t�����'���9:�t���r7ѰQ֬�Z���C�&��	��*u���m����Pķ%�=0�3�K��U�#�^^nj
�u�Y�ee�F_b�����$�y��V�A��4ڟ���Θ޵#Ugvv��}�C�D:���S��ל��:�M�¤stI�bV�mɧ��sE4K�'.��'u6�����t�`Ϋ���.�������p=a���y���3RF5�xxڛ�j�X���yE���C}T�\[������|���]�U�p�Ia�1����~�V:惌%E����	j��f�.����ub?���p���%S r��������*+m�kAib��V�f�?O~q����f��F�<L�qo8�R�j��}��n�w8������բI�������J��V>	j4�UV_�C����0�\m��a��'.��21�?mZU#��Ѽ��@�@���؀�=�MO�l��.�3"����n���M�T���ʒrg�q&o{�g�rc��@v:�d�:����D��h#Gj=�e��o����͓<��{���'�~0���f�0���=�Φ���Ŷ3�ʋ��g�>�dW=����/U��I�td�������'��c�:�9�F����=aWOK�&7���Du��Z6��I���az����b���p��gO��	��3@�b(۽v�ܮ�മ��i("ϟ��d�詑}5.���L문Z��l{[c{����l�E������(��&H�����z�rZ�d+fdI���b6S<N�J�����m���n��d��j���)� 
m�Rr�ᢱ�a<.u�4�g�O|,�I�Ȩ����s�څ�㦗9�SX��5�~�5�}�jD�j�
�l�g�n%ݹa�pgV�/ۤob+�g <���� DѫI.�JGA|S@w�-����B|��߭����:<�M�/�/y��*��^���v|ZY���2W������wS����m�
�R�턎 ���l?�����]���~#��hE@;H�1�.�>�g]h7���W܈l�D���|>�ue��x������3F�������#!t��}��8ɑQG%n/�-rWz�´c)˹m2�8��b�����6W+������7�C��o��)���o���. ��eY�Z���L鈙�T�bfoN�	���1|���*#8s�8�ڙ���Rŝ��
�9s_�H76U���~��A��lNrԜ@���u�L�R �[`����8�iB�{4T 2ʱ�uz����+�U��=�Y >|����t���H��_��H��r��m�f1��TVom^���S]�W�=�.~~s�V�Qp�S�� q7��ȗG$��t�?d��·,޿�6�RP�|�;�'0p{2�����	K].U��|��HQ�q�-2��>R����!֬w���jDQpK-��a�?�ڶQ��Ԕ�$|7��)xPO���3<=cs>�A����Ħ�	@/��/�'�k!��`�=�/�g��b�E�p���	3ϑ�^�ř|�(ȑ�2B�8``��!�U�n���E&�~�fw�	Z�(?��9���Q~WVhkFS��F<{�	�H8� ��d�ȣ�8�=1зB��Іg�7�%��A�ԗ�m=��Jcn�2p�ƣq�jD�7�,*�IC�5d.|^�X)8�<��#��i� ���y����؞�kE���*��Mp 8�5�޺����eGؙ/[���`< m�)��[�����y7�����I���>"ikTe�����ǌ�H�[��#�(�Ao����X-�n3eF !�B�J��_�g�pj>���ȍD4XU�����Jԭ[e��v ��_^��i꥞��& �l��i��z5�������Ol!g
ړ�R���z��2��3p�@��/	�;��9ah�wG�0������$
&��мPۺ�²5��_U{�S�k�f���V!@��rd�vиCW=�SBXwO�[l�<���Ɩ7���q����Z%a�o6����$���7���ۼ���������]����ނ<�i�@�#���Y��u�0�`"�K�]�����݂5�T����CWX��ٲ�ó�V�,���_��|�����Y��IƎ\YDś4�(��P pl ��Қ�\H]�wS%���A-�G,�_Zj�t�7�H��>*��0�-��2b)-��/x���ިS�=,�w�=:Ń��d�* H��ؠU�W�7;����D�Y���]	[T�B��ۥ�fS��8Z��D�v���J�j�_m�^�挈��*�Q��՗;B�i�]�ԊQU4���È�l�	IG�ą��w���P̀X����FKdmx�m\��!֍7�,�}g���� W{��=����j��u,�,h.D��������x/���f^8(,�6�p�B1�}�>���
e����|�C��:?�j��F~����n�u?��ϨƼ��'��#�/]���%\YU��@��8e���z���'R.�ླ���g��xl�Y�q7k{����@�,|���O[/���w��m@/r~B�������O�kTZ��b�>�(FW�<�"��k�$5��uP~Ųoa �[��z���ހ���zH����iJ
�@n��R�-�{���y5�$���i�Yp�l�	I�c�? �	ɀ�uh�)�u�><�BA�S?mW ɴ�sP���R��Nh�$���R��CP��-�J�j<C���2��#5��9��~�����]�?���o~PmE��N�D����غ���.��Y"=���W����%׈�~+{2N��ڍ�:���j8����ʹ�B�X�c`���4 Ĉ�NW�~� ��)f�b�ԩe�d9s:W4����;�݊Uc�S#�� Nwwg�I'�ˮ�Km�����5z,�S��Q���5P��}��:���2���,@6�{>�	 76�d�$�0z����st`|��D��}���h��c�u��'������T�20��%<l�t^�h�{�lkn->|��D�,�q,/l�Hgv�?D���A17�����'N^���Jik'�=�Aj��\w�&��w%B/^�$0�a�����A|�
��H|��+�1?U�gS�qޚ��������'�2<@�'[*1��Z_qt�=�tC�U�U������ ��H��[2���ݿO�p *�'��sa8o�>���Uu�)H"/cwMJ�x�q����^�#�4x���'�JN��ާ�yuwxy{px�EiNH�HQ����0;�e�Έ���q�\\ΐ�]��9蠂�El�������S��?Y�뉩Q4'o�<�����e
U�݋�[��S@����;�&�LL�	=YJ��BcO��ҙ`�<�4��P&�:n��\��-��6����>����K��щC���:�CS�=f��f��\�'����U����f�EZ9��S�:t���1C�NTѯ5��/!=Ib�`Kŀ����ґ�_¢Xd�M��K��yL��+� 9El֎��S���;�[Ӹ��Rn�˃GtT�����p�pq��k�:�7>@#\�'�G��mֱ<,�p&���o������ 4�ӽp,���BUڊy���˘�"�V$|\�9|2r�g\�;�<�(�L\*�!?E�K,��{f��̦q}O��X�=�p�|���r~���_�����Ub��z+΁�%o�Ti�ndG�x����V0�W.4&���=1���  ���=����Hn�5ޛ�_TV�g��� �͓S��>�A��d&��C���Pb���6}7�n�P8@��\4]Y%d܁|�T��-�&�ԋ���)��y���w��V!��Q߆(Q<�m�м�M�5�"\�R ��&^�Nge�΅��5T@���.��
L�B���aYK���w?���b��	{���*Ӎ]DZBӵ�������\����8��b�:_n��4�전��������()X0GF�۱����{�f��C?f����A�E�"� 	�-5�6�u���OfMJ��6�#� �9ʖO�t�I��8OE�gH�ݠ�j7O���F6�ۻ:�o�^қR!@@_ycVf��ΙyVk��=f
�]��)�.Tޖ�I���4	�;io��]�T�S1h�.��l�C� �(�uq	7�
.�<�|ܲe|���?�`ː>�E�vw*KO��pOv}����	k�Ue9eW_1���k��"�]l��D�H�7p
�ɀOiO�W�?Wh̗����E�"L=̐���I�_�g���/�ku�R�qi�|A�lH����@��ޠ�&|y�Z5���6P��*�a�JcX9�2��Rf����D��=M�C>K�8:�x[����1#^���mu�oX
����?qTfI�o\�7���N>G$��Ť\o��H�8XH��5.	g�a�KC3�M�k���ƶq��,���X���-TG����OS'[��� �h��]�� �˘�!����4~`24���sĲ��vx8)�^�A�B��P�ǗF���AZ
��rOt�P�X7��3u5���b߁,�e��_�kt�0��B_��" �-�s���N����n&�(�:�dꮯ��`ކ}�_��lВ��	�t�2�0"���������Wp��$$������<��<�7�( �=9����3�+;�����C����bK���J�kg!�����)z�rqܴ���	��N�Bl,���dp��c��kkA��щ
��6R#muny�+��o��W�S��q�pJp��Q��OD*K,!���u� �g�{�o���o%�ɺ}B���o>���^���F���~���{�I��<KK/￦����`v�]�8U��a���&����Y����-�;�\^kѕ�5��gm
�:m��{"�r�lצ�x8���&5����1�,�J�M %��í��e�,���CC��*�^a�Cl��[��)�$ަ-��`� /�!z�?Eޯ�p�)2�xR�]T�\�� ��d��W�����q~���c*���rh����k+A�YY/��ѽhr��3š�H�z�gm7���L���_��
E��u�����|g�y>��KK�!\-�0�����կ���8�.�y��
��o��h,����fUԀ.[��/6�z|��`V��8�B�t/�7 L1;F�Ԉ��]�m��T;���/�l�e�|ZX�S	
c�4���kt�v�T��N��˾�����W�{;�6~bs����e��dx&"��k��w4�?jV+���y�U�Nr@����!�h��`K�q��֯C�+(̶q��f�M�m3�һ1�(6��KcĒl�e�n��u"̼O8��� �v�b%���P����k}�);w�qP�<m��{�W��ս~vf2�J0NX$N�����]0A�n�85��w��*F.Dm�zA�e�{	� ��Le�9'��H���Up|����\��mJ��3��
�#`�M�zoB��zgw��-
�`.c��q��H�'&�.F����ЊpO��?��N���J����
s��z�*2�Q��hn��ǖ������wi)�6�
5������V���єS��4��<���?����KC����M�&��[������<fڥ��k<�����W�&'X��3�eC�K���epj��դm.U����N[׺l���c�'�3�C���F�ۄw��@>:�� b���/��ع�D���� <���R1���7�H�T�1}�e�����.�#?
l�Y�Z�&�X��V#p�Rzh8��m����y3�Wk͑�۳Ϳ�X�i���\�S0&��Dʠ1!�.6�ҽĮ �F+���؛n�0X�_v��82o\3t��0z߫�����aC�͢*���_��J��>vح�[B�J#D�)_6�8z�'�o����l-�*P_�(��|����O_yl~�b�j�p���s)�<�Y����z���-���	��J�i�y4���*�%���	(S�?���j�7(́����1�ڂ�נXBI�ڝ��-�)D?R!v5��7�ٌ����/�޵��ΞIP�h/��Z7�ml����%NB�mZ�#x�8�5���4�� �i!��g"�O��퓷�&�ͤ��_üU]L����b"��-Ŷ߄M��m�y����&i��r���ϰ�9�װ�|;L���q����W�3ZL
�\�S+T�M�<`m�f�AP,�4��7��eB%@v������k0w�������ϑ��l'4g�)�L�v��@���'����>P�Y�nZ-�=QCǼab�9{3�.ˋ��	ŵ2�I���YO@����xg��S߭ٸ{gEm+�$}I`��E���������[�.&�?���C��W�2���Y�h�3Q����v�ͦ���̚�\5;�s�����U��`��iȑ�a�̯�N�3 ��,g�#�a �U���6�p���}7u�6cի��{��!�lAv�CM�_�kt����Tˤ����4=w:GN�C(���������9>�*��WC�
��v4��L�-�U�����v��)C�TY��4��)N��8�\��yf��a�������l�;O�β&:Q���7��w���[�3�'�����Fr�7JJ�i�t��e��z���� L�u�����oKݻ���%ر."j����q��5�B�5�������=Ie�?�p��)~WDI8^ѭ ��!�������BxJM�o���A��o{<�W[��.�w!IX�������fW5H�z��x�<�!tʝ�F=e:�\�/[B���L��y䁂�R�#�oG(���L|I��ĥ�x�b7��K+�S8�C�T� $^���6�'=�����ì���������P�e�y����1X��8����̒m�e!C�/|=L0j��l�ܾ�X�ȫu�	W��z����/�g�9|$�����j��3nˁ=��q�κR��m�� �������:dr_��*���|i�{2`���
�~�NG_�rM�r>%w��$�ʊ峳m�ݯk��#̞��<����'}�lv�g�^|�}˾w���9�e�w7��}�fZL;G��A��ZY/.��M���g	z����3��s��Ճ�����W����R�Y|j?}{hc,돞�p�9�d�>|)+�@|��;;~�̽l��]�tzk���������ΰ
GL��(.z;�_�C�H�{;��<s���F�D�}��x�5|Z���6@h��c8��{��b��}���c�t��IV�+�����p���[�8`<?:���l3��J��������7�� fcx��U*R���˺���/����^47��)���'�.��c��t�\�W�	%���u��@���� +J�u��.�y=��[TdtFJ�X������\�����7X���%"ӏ ��M�Ff�%l�
��r�l:� ����������{�8�;Z����9�;�5�s����*y.��q�-0FH����x-�%��S_�`s�?
G�l�/m��¦�q�(F�0yzZB(���ƄKQĭ-��;7�</ۃVg����CC�M2W?:E�۶��^���jM)���gOٺ���!�\d�^�����!�7�돟R�����V��ww�+��r��r�s]SV����!��:5n�_�������>��b��t��[j��ϗ�������F�~B�s���	j$��_;~<���c�?�FC���h^����(�N�.������ ,�7�S4o�s��/liO��a�W	�Q��s��x���8�@YX�ڌ���5×�͟����g&)�(�dzUz�����֙B���w~�	PJ��(��R�/�а��%����uv穸A0���U����#8ӗ�ޒ�w.ԟf`�H�'�_@��2��č������ֽ���������WY_��mz�!��%o���m;3-t���A�����.ի�u'2<�`��'t��;����kV�;��؏o������������J�L�G.τ���Q�C�߃������%�Cl���7����(��y�̄��O�W���!����?vNR����Ք�~��è��Z�y���[Me��5{��a��l�G�T'N�����,����S�|�?LM?q�M��	�.9�+q�����ލ:��L'#�s�����?lu���':Vx���\wg�?��S��Wo�i��?�;%���j�o��ƞſ�ck�t��o�������o�ǟ:����6Z���B�o������%E���vY��4h�S�S�B��尕���;�縼���c�ϸ/�i`�}�?��@,��k��w@�ے.ʩ?$�X��Nor(;��������r�2@)ALh�C��V|e�`o/J�e2��xye)3>�>��cs���P����JPZ��>�%��V�F=�r�^���Ə����!�яr-Ƚ���ƥ���l�����������yyҞ�k" ��"�Y�\N� �/�~�1��!�\I�/�x��z���u(SX̪���n���5�p�R¡�2C�o���{mscv��;��ީg��VgL��=�[��1�v�>���Y����x�I���N�������$��:u*q����&+k��!���Y�qQ���<Z��4tc�_˰�(��x�z���2.O4$5�CR9�%m43�I��2��κ�&�&�rp7S���ѣ`ܻO݉�z�]�fl*F����z6�g�/Z��c9��de�"�;���y37�c!^\&3�|�IE���l�/5��j��D����2ֳ#B������9 ;˙�ǬWĽ����8A��u�2׾�j&�K���b��јuR��V��%��UpKB�G"�Uvm��Xr�i����zx�)�_��X|���zU�3)��=x�RB���G�OuMc�V�Ē�fp�FM��G��$'AnM����U�(��m���?;7]�0�q)���\UvQO{����pQDNN΢��!�����?K�l_��Ai��O������L�U���z�ҌF{ٌv\|(�ט��s��g��82Z�_��ik1�R�u����lI�#/' I������N7.�=��OO��̒u8B�&�x�JT�:���bM���j1���g�xO�ȃN��_� Bm���)���'	�^v,u6c�j8�K�lp�=�p�y��̮Ϻ�n�)��P"�*fx�������w��ߙCG}���vkN�~���C=`���_\t˕�*��s�z��UF®�/�~8��i�i-�3��+X�Ց�XQS���_t1���J�k��J���C6m@q���E�'��h�+`��̙m�/����q��۾y}����Q���@#�2�]!�C��I|W���Z�����֋��*��Xf��3����	��w������HX��s�Y�5 B�N�Ƀ~q >%:<>���~���V�Ǳ3uL5���� Y�*]�?��4���Ξs;���~���S��ʷ@T�%�]��_�� �8����6 6Q�f�YQ;��[�����3n/���4P6�,���k$LXXP�KO�zWs����ܻi���W��d+=�i'�B�x�}��M�q�V>�u���ad������g*�?���z2x��3�Ý؁�T+SS�c��xA�$e�zs#�N�Sʕ�C��E&�n�Zb��]>:l�w��u6����������b�Ȁ��,���ݾ���#jւg�۬H���>� ���v���X[�B�?�qq���8���g�J���~| ��շS�1�~ޑW�H��s�m����lVׁ����������2�J%���-x�=��72�&ZV����	�*�d܀��i�܈���� #z�W��|���_��>{�&B՛�.��p�����e70���9Nz�}�l�s�?�c;*_*�Z��/p��F\���6|��L��j�n�����R__�M�9���=�"e ������ ����'EF�y7�R��א���6�j����X<kC��(59S/V�����w"�U��6�'���*ڃ�×��8,G¸�
,�s6��^�>�r �캦�E�Z3�d�y����0R�����(躴���.�r�[ oiK<��W8?�j���5Z��XE�5y)敊�����
�%�@'�O��u40���S��wӇf��K �4ޞN���$X�2Q�
V���D�~� ��dM��%�V^Or�o3�6(�3t;14]=�����>�� W1u����Gw���?gi&�օ+�0g~]��O�_>���������c��XU�T�q�G�q��aI�ugF����b�ԬdpW�7fr,~�[Z�ߨέ��΂|�,%�S������/�g�{���8�n*��ӿ����3�N��Gg����_l�rJ_��f�������3h�t����n~�I���>[~����G�7� ��sF�3���0�#e��^����>ʳ�HWO��k��+�TI������iަ#G�!�n�>3356��H�!ӿ	֊~��J\����Ј�S1���	Ϗ`"m�1+��P��� ��:�
\�?��U.=U#�ap�[Y����F:L�]`�,�陘3���sw'+k���L;NN^�=ï(�c��ϊJCi�(`-�	�a�S]Q�r��o����74d׾��C�U*�L�H�

�JJ�����l��_&�cq�p ɲA�!��i���!צ�n��"�y�ǃUh�[-@݁4 �kbr�`�Q�
�68h��Zp���d�!�Ax�
�>0��G��n����ҺZ�P�h4��h��E.� Q��g��3N�w�v>�����:��j[&X��'X�_�1{�yY$vƅ�1�[���o�F�~0^������4�5�'�j�u��x�O#�ѧR%mF���߸_�A����Nn�qvYوG�@M����U�IH|yي�nO
|Oz�DD��Z��z[�!m�����6��
޺T����RP��"URlh��a�
��s�U�J㺦��R�GՒ��Ao`l6��#�ܜnXw;"�ײ+jU��ƽ,3�=P����{p�8��˩���ӛs�>��q��RD��VH�Sa8��|ܠd�"�k9����T�IQw[�����#_e��+��*�n�����)D�T���4R)|ʞ�'�I�.xۼD��.�D��:?=!�롔fD���P"zt��{L"�z���ݿ�r�	<!�ܸ�G�6�V4�o]F�t
�t�|>by�w7@.�L�b���xvfR��>�ΰ��]���S��4ڮ�Ũ
�ܕȩ�򜟁m �9�;K�2a�}��܀�XY�觑�E0hb�^�I�t��m��w���
�h�}8��=�@�9�@�z�-�N��`��}hN�_��ū��� ��T8�n�9��&y�x��8����|�r��4K��*�)Td�IwWX�MPRJ�HUѬj�i�M�a��]��K}�c���M!P�;
a����8-���p����Ր_��apj��ኬ�r(<1 �7�YY��q9�:�2��Wk�s��&�.��ˀ��y��Uy}�C���r�B2Oi�j#=2���0�~dT#hw��a:�+/�u͢���c�:��/YaQ�[�F9�
:������o�\��R�J�_��x!J��v�� �ߋ�E�D�����} ���ű�>-<w��E����Q$����,�A*�X][gn��� ���;
꣺������הtP]��\�}��Aq�2P�/�(Fs@kPfo�ݹ��Qhk*��k���;�}�ړj�5�������V��N�޽�%����\�5aeӎ5�S�+O�PS���=VE	{��+%OT��WД₁��i��N(�_���8auq�P7���K*��Bؘ5C�Y1|�j�J0�pCJ:��]*��j�l���̏�${�h��#_sk��str1�3����a�b�	��5{xlu�M<�nY��k��[�mʭ�?���<6n!�Sep�,KX0�wMM �tK5:��	=d?��8�x�A6��� �Q��� �����q��	5������R���+��r�H����<vA�aXM�hg�p���	.�m�x���	9 BYywV�����9����8&����RR�Lg��)nQA~�i�u�q����H4�M^���>)���%�A�m���q���z#�����}�ŷ[��)���N�>�l_7͵�c���Y�`��kA]����B�A��k�����<r�_ǫ�����YKw|ނM�F/�H�����̓`�9�Y����)I� 5����?��o̙��3�!�y��ׁݫj.q�+����V���4z�cn�x�Ѣ��cg �Jg<��j�jY\'b���
E3.����1ax�D:~��ky�G��))����F����e��,�m�SQج�K��V_�#�ou��Q�io=�e��|~']n$��ѫ���^'�`���TA��)���z|�x���Y�aǸ�R鳌y��c�_����pfx�$W������7��-��'Ht�6�!�I�^3�����#��K��}
i�8�T�]<����j����N!����|�?}s��v�����sۅ�A��qYvݛh9x[Xc�����ַK��!�hh��<90����=�lV��ԩ��ޒ��0��ҽ���,��\�F��7}?���ҽM�Xb�m��Ì `Ð�o{
`���{�Ǣ���9G'�3�����:����#.s��3���:��3u�!�:���o�B���ɋ���-ąs}+e�����5�mx��I"]���V�P�ж��ï��痲^��k���|Z�h�I�2*ngXTU��F�nπ���Q�C�|7�Y����-	�M��}m��T�dT���<��q~>Z�
m[GN��G@�yw����u1���df��f0�{MM��y Nd�(�f��o��6
��l�1Q�q���H�Q�c9�m�D���ʞ�i��g���٪��]l��_V���D�C����)�A��U_ԭF/f���2T�)e^�"]Ykj*�(�}U�s��^��&,zX=��v�C�x,��%��ILqJ�c"��3����
"�(1޸�hv!	%�P 8��b���KĞ��o�I	m�'G�<G�mv���`�~�R��jF��}��?×:@x���m�2�6ǉ�\�ܜy��c�D�C�\���pg���M��*���z}���Z�PB������Z����`��p)��"�N��h��B0+�"�n��\s���g�5��_opH@�\*�1��������p���;�nŜ0^�N����2��8���'4��wMLOsW�r�WW���2v�N��ޫ���UupZY�� ٿ�#ML��>���&�"��a��kP��-𥑾Г�߻_��a�7����#�'�ݖ*�٤Dt<�7�0o�����㆝��!#4��_qܫ8����Fb2�(�+�_��	)�Q]�7�nr.*獌��M@8�|38z�E\���g^�zp�th�+<Ae�?�k�䥾�UΠ�8��#�_L�8@�mi���±��Q���+�us"Zi�6��rT��)q�%6�-���E�7����C���@�J��͂͞����<G^�^�A��P�Fɰ회��Oo`e�m)gC��"`ogl�<�p�-�0bfwabxأ/�c��RA4h^��݅
����%/��m��K7aJ����{S�D�~p��a�ڣ>Ћ������`b�!斦���v����5����h�S߭7������F�A����FWö�u�*B�^+?�Z�O0|I�F�[�˺c9y��_�i���=�P��k�ǎY���N[M��w�dO�h.�	�:Ǜ�Mq�
[��7iD��}���?�7,�NQ,���85ʹ�U.�@�q�-��J������J�/u�����cGN
���D I�	�B!o��|����~�Y���6 ��;��#|��b��ZP۬�0W5{��f�7y\3�p]+�t��p����#�����/�,�*R�0@� y����Zv��[�O�::���*4E���꾟U��\pF��@�'�b�Ar�*%��5o 3�/-o���d5�x
���r^���DNJ](�Ky���j霡i9�e]X}0d�|�`aN��L�B)O@���˂X�"eG�`�Y���0l���e��v%��[�����}�>��ޯ�	���1fD� ��zĀN�L�օ����
���4���k^���i�d6S��������?�6^
��
j+BN{85�Q6�^}Z*�ř�fj��F3�G�<mC�=�#i�ݠ�h�_�<s�7�{�~�� ��J�K��.��FD�c������O �:����QXI�]��pϧ�'rrj�U�K� ͳ%])h 40p�tV���hܜ����h���"�H�i[B5k*�]g��dӪ�ΝeW��A�Y噭ݵ��V9;��7|�A©R y�eWĂ�5ս��ƕ�C�����[�Z$B�BQ�d�K��!d/B���r��>ٳ'!Y&����a�-�`��/����N���ԿO>����<����93��.�ɭ~3���+��J]�{�R(�iń�w�1PEnrvW�y�������E0� Y�n�[�M����~_j�#��{G�w�������W��0����%�G��s�ژ��S��:D�"�\���	�ť�*M�n~��2g�v�O����3��lDҊم,G��G�v��/�n^F�>�8�z�-�?x�)(0]$|�(�0Y��|���Y��^nwi=r���ȺC�*���AAX4�`en~�3n7WZ�ѻ��S�2��<�-����%�3ښT��:ZL`[N�~~Ym@����i�e�b�!��f6�h�]��|a��Φ����������Ja��a���en\�]��L7������(n�&�C6�b�{�e!���~��_��4n�U�w"�F�r x�X���F���-V�Ü4�R �v?��9l����׭�*�8C٫��}K0%�j�����Z�)�a�ʆ�qȍ���N���:���x�^%�0g�f��lM,���n��r&~pF�q�kx���(��v�	� �����kRȡ=��VU&o��z�!������~����'���Pb�8�?_7�%��7	U�����ٴ/��F~z�@��#���풿�"GmN-ڡP%.�`r�����ps�������rٟ�Mnr��հyU���\��Sޛ�A�,���2�S�K7|��|�E|�}"m�)�X`�M%�r��G6��r���v�:!�Wl}����ʦ��#@8t^�җ@����'E�q\Z��5��)04��g8�`�]w������y
S��l��dR;iJj_{���+:�ѯm�! rK�n�r�2xct{�`<�# o������}�=��?*@�����!oNZǄl�u��}ʫ͖�'�6ޱ��d�M��d���y���7�Y�ٶ����g\nX��7����?���BX�&lgr��4,�L>[8D����=z�w������^!�D��2�`#���ڱ8��	�)n�'�LP��6K�@2"��@`rȖ�B�����!�h%�彰�3|����R8E�ƽP??����btu��[�jJ�4G��U������%{ԭ��r��Ȏ�7ѯ�ܜ�/x�[��v3'���c�wK�W�����&�d��b���eO��^���̆h�!�n�n`�&[~+�4!�ޫ���ua�ެf<ٔ7$�!��ng�B�����~�n�y�@E9��P��1���Æu�ס<�PJ��S�71�t�l��B�}$j1�,�VD��F)�݂Qo�=���c	�U����G.���ʀ�# ��":� ���T�F�߈�y���O8���ޘ��T<���4'5�sn�K���+����l����|�w���ʤ�
�Mj�c���G2ɛ���8�d�L$G�F��5�&��/9��rN�}�Sj]�B��s�V���n��x���U������񻟕Ad�8����o������S@;�pD_�4�j�Z�Vj�ǃ;�D�\�����VM��w�٠}q�7�k�mk=��u�K������~X�}�����n��{g7�?0��z�}�8��>�M�kX%���ū4�>�K"�DF�ȇr����S �\t����R���]�m�����i��d),W�2G�c0P?tw��T�6F+��B�^;�R5��[9g����D�(6do��-ph���e>u'}T��ܕ�2S�cC]J��'э�{ۂ7J`P7$��Х�D�屌TH�"�(n��Wf5���=�	�i���Ԭ|�q�'_���o(�#�[����)!�c���#Ĥ�Sq?*gBa�ȡ���`�޶�-_y�:����]j�ZG
 >���>�f R#uDB|��ϕ m�1���0.~ ��ۭ&PT��qGȭ_N�L&��)m��E����V�^��W�:�/#M���i�S�����������Б�q1@9�K=�?�F�Xg�/�d�y���K�.��y/����u0���.H1�8Ҹ�*���+���w
V��ծ_�x��UG�U)r�Rt��K��	�n�7�L�{��+���mr�#Ǡ~����v�ꎡHSb�ru@������v)m�m�M깘
֏��:,.�LRJu��cR^���|8���)�3�1~�Ȋ��3?؋��oUN&�����u-��#�F|�*zS��I���;eH�ݠ�5ٸar��*ò��.��;	>Ə7�Ef"]f$no��޻���K��sy���	h{����tF�yn�y7X���J�O"�������j!��߸ힸ���9Q�Ys��dse���70���M�x^�2� ���A�p%���*��N���X;ĳ�D)?��G<IѠ�ć���Y���Z߬�Ӱv�8Z,\��3���翕�t�?^�J�=��Z�?d
�����}|-�A�'j:�.��W��w��Ӻ!�_�68��\�o�JE����/�a"�i�?��ݴ���g��|s�����@_Z�_y;�+=��?��� �#��x�^OP�DK�������hU����_D�	7{�����2�b��L$��yՄ7�����&n�ާ����Zݒ{�k�?:��#-�����֟N�y[���ҲmIwP� ���t��o�Xs��ɂ�妁œߩV����7q`kk�Z��p���K�b����l77�/�ǵ�;fb��dI���������ԯ�L�-ˌ��[n��~k�ﻥ,�#�׃�k���8ё����*/��҆�9��\�l��	���{Z�B���h�F��}自sW�Ec��
��?-���8�N��!�5J�J���I �3F�g�0���*�������!��j��~�9L�.E�&��� ]�W|��p��~�}6�`�H��gG���w������<W��N}�,2RUXc���:F)�*%��E��|.rs��F�^Q5�W-<����,Cۼ�Vmĭ]p��{~��zc�� Qo��ǈ���;u��9�i4%� ��:0JV���6�
j�^)n�q�����Z0+�cS��mUiu�avp���H�<3�N�6��{bY��EQ��Bq�7�[O�4�:�Q�g��z�.�q�,��-.r�<��ءW�]~�0�YM��P���8@U�s��C5�w��Wk�5�:���,C��,n2+a�����dz}OP��n�&��Q��
o��qY3)��F�
�:�F|�S�w*�S���v�@jKy{WS_��wd�#wT������̟�%�uA=��#kU�`���bg�� �����0��F���;]�bb"�-��O*EtKy��9�߳J�
�� �����KɅ��u���y_����="�fs)�0������O���W��ǲ�X�bL���Ji1C�ǁ��Ll}�YSl\�d�*|��rT=t��ǿq#wﬆx��x/oZG��`���йn��$�
��7}{t�dl�𰦶�,G�C���hDh��m[�c��z?��@����������o:����{$��H���x��j �8*"�֡���R��3(��6��D�&e�lX�����'l)}N�WD-�":'y;�S���r �i@S�9J��	���sYŨڋb'D�gl��+��F�'�B=n1%���_\�S�9C�۲Wh9ejU�Ҿh3`�H�ܴ��O�l���1?�2��^��y��b��x^��&w^��M~ػ:�(-�uSh� �D�=K��0-S�o ��n���ρ�&)*�d��EV�OG�+8:�¥�H���S�'=�υ9�=4�h���~��T���)jB��).+��l��&�ZDx�"�J��͠mӥ0���c:�w#>c8�!�~�p�X������؏dq&��hM���y�3a�3��ZbN�y�b��uZ3��������+|.�&��F��*�uzJN\3��S�g��dH�&�rH���އG����Yv��\ΑU���^���܂P��ɦ9dP�e�8���;ݟL��[��G��1���&�ӷO���sy�������Y� }UW�9]�ï�3��H~0�����x%���"ȽF�I�<7�V�=O�އ��p68X�j�,��D�"Vsp�#ܩ�;�޸ی'vE��i&s��Y�*�1&LN�o��d�,XWO�ڭ�Mm+2�R�̙Q~�XO���xp�D�"$D�4v���Vݠ���ɥ�P`9�����iM?��m�<���D�\0�k\�2�d��U)y�/
�-��(پ-(h��هw�c�:��q��aQ�y,{�P�^����E\#�� :��w��:�Θu���AK;�*�2C�ɞ>�[�4I[� ���W]���"��v,��0QA���ތ ��h�[K�~tY��wa�u�n�5�Zz�b��-�3���%�,h옐�ps/�K-mfs5�,bl���Tbl�-..m�U�S�Mŭ��_ki�',������=eY; �s���Nb&��@��ŋ7����r��0S�w,���ut_Tq��	�n��]A����$;ЇG�^i��G�<~���2�)^,�-O$�Y\�+�:�H�U��}�����D�&��F����Iu����9�����j��-W��Ś8�p4�t,�[� =A?r%x�w�M�7kfq�U�B���$��L�y���LM-��Hz2��ꨡB���3 O�tfS�xyK��)�����6��oK���Y\}$��z���aϪ�!{VK@&0�۵+���	�Y��WO�K7��EQ�&v��Ҍ xF��ۯ�y�}�0٬��m^�yQӪ��.*+ˈ�  3a���<�R�ybT[���Y�?U��ҟBr�@�j
����vN�	��{8���l|=.E��d?F�������w
ao��@Zo�k/{�f�шO'*"=N�Dh�%6K ��)���i"�鎷�Y<�,���
mAV����kW
���ptYw��|����O�B�cJ���^�����		drB+�H bu���/�	T�j�J6�|�ؔ1�a�[�x.����[W��8�<���+�ezMg�,��BB e��b�U(�q���֯,�"R%m<mT�Yb(݇l�}Op�-Su�cbӒL��TֳZ�oZ�P��Z;�$e2'E��ج��(�uO������r<q�;���{;5��h�r��p�i�S��m�`�Ym���lkc9��:�
#kЧ��֣2�Jkp�Ē�(|�ئ�X%��`�T����a�%0�P�EUˀn>��ԟ�R�ý�U(`b����]ѭ-b�YhkE��_p��`�������]�g��(kT[�=SӨ��.T�?Q������� @6��U �b`e.�<�����Ll���0[C1��;d��bn�<�z~�4 �ѤV���/�n.OV���vy���Rr�ܞ���Ad,H�W�P�Y��T[��Yc�p涎��K��rQ�׳N���:�<��?2y��=���<H[=����H��UO�^5�pLML.�nS^,��&��K�mV�Z	P��Hf$��.�4����ݛ}�6E]��s�G�$O�>�.��z���v���j"���З$B-��-*/)����ѣ�}��Ԫ��:�~=Pj���A��u�_݈�q�� bXOy��=�V+-1R�_��s�2�LRp���)��V�B�:�{�H��η)�n,j���GnU� p�U�60Y��Y��	Yѱ��.�Vӏ��,�*u�z`��2�(��y,�b]M+�l��m����m"}�o˯}���7#059�S��O�(^G��[6��7Cu��pu�;��%!��X$�C�G�������F��j�U�����ZN�&������)L�R`AЩ���Ԏ���3ۿ�՜��Ď.c��(((�#�Ap�aZ�D�A��6[8 �r|,ܙ�9�`~0��B�-,�CH��Օ-�&/�Y���J^f���e����/��#nQ���'ϡm_��;�.��l���<� ��/FM�ǻD�$\����1�^,�S\��=D�׬s����x��c���2��x{���r�m�r�&�Tsĺ���$�N5����\+W��S���ۇҤ|�7%!ءG��/��S�]��]\��_�˰��8p$ӫm*��V�I��I��q�QZ1�m]\.2�(1�E1�s�`�w(�� �P��:��:�Yffy�,�=�n�����߇���^I*rv�����qU�xQ�;���M��+�h	��id�}dw�m�%ȍE����(���>d�h�ҁ9cv=��M�u���L{�AB�����JS+����v��wb��߫H�����_y�����������{���6��*�Q�֍���:��2=tBTB�����S�k+�Af��ؤ������K^��&�e�U,�yn�[՜;����6�3���~8�����/^�t��=�1j��x���V�N��ej�xU��V͢���¿=X����U�]̮&��h��v�+'}��y�j�adahh�_b���vWD=MR��Ir�����rD�m�t�'▟*��ז��^SW���b��i���vwwKIb"Y
\--.�f�6@�V�	~p�K��ɍ~����slur_,o�d��%����*��S�k�mш ���l�6]�e�g�b�9��X�Z#�Í���A�+��m�8�5؄�3��Ok���E'�h��Fa��,�C�W�kgIt��^'6��F��喥m��>��� [�u������XRLL�q�le�;w�!�'���.���I���A1����i1�-�;�
~<f�X�����c���[*�ҷPA ���x�;~)�I��Ol�����T�>�٦$P&��j��#�#P/�_4zvW�S:}�j�O}�p��Lm��+��]���]J��'7�s�<�p��q���_J�u;��V�F��
��/}YN�1OJG	��a����`��T�(�Ԍ��3 ��'O%���~�xFC1<V�' .D�JwD�
=��I�V�N�Z������e�Ԝ�É&Cz� �[e�fP^�� �lgj�	�ð��&�k7T-j+y�����JK�<'�~�2r꟝6����唭������U����c�{�a,�r�d�pс�G���I����=���2<!*:�1�0�{uZ��D"w���N{��4��t�!�O�"{��h�=�qQ��8<l#;���5������c6��:�6
9�@��,��˯�㳐��c��!�K��@�b��6C�7h���(ZO�̬�4+�Y����e�Ӻ�����'}~+��}ɯ���c��N��g?=�~�~丰�<:<��2sc�Tˠ�����U{gqK�C���)�-�Wj!n�WX��-,��I��<�bq�4�R�y��,�;��x��e���J����s��zG��{��cn�����#�5q�&zڱ��J8S�dK��D�,6Z��խ�F��~��zΣ��j��m�j_o�D7��W+P`>��Դ��oև�]�:m���%n�/�0�+����D�˜�s76�I/P�E�Jt�I���.un��\
t
��풆�C@�Bgj�i�D�V#F�9,�J�]F�Cگ��Q������'*P�uA�i1%*b��VO��^���8YS��Ѣ�_1⊄��kmHn���j�����f�YP��՛,ΙY2G�����y�.���Ȁ�{����/Y�"lrns]"���<]U��9(�u��*��}����م�2i�%;�-L�e],����3O3Fn��;��q�^��M�ӊ��☕���րe�3$t[�VnJw�I �C����i��s5D瞧�G����4��9x5���7�Qg5v�@I&&���ol�Ah���Q�CV ��o7�mҝDN�eKT�c߂��}�P���	Q)�L>jmoH#��.WzV�AS�w�&���cN��07ݖ�G�lT+�0!YPzV�ֲڀ��Z��l��.��d�������x5jIh��QIr�gI�����ˈO(B�I�7jjp��w.��w�yP3IZ�¾TR\R {��P�ݩ� 9�x^Q�R�0{M�8���t�b8n!����q�]QX/�1���&#���F�i|����,
+��OI/yip��>0��8#��<��g X�"�$ިЏ��E�(Vc���{tߐb1��ZD�9���gW�(�1h�*_�X/�Dm֫'-Da ��t&��=�<��{��$��@?i3	#�]SbP���|g0�oˣ��-�kj�ai�9��j
mY��
��[��E���/K����!TfL�D�b�eccUB@"�F4TGM�yW�}�eϮ2] �V��<u�I�V�3~�W/�\.o��tAL�qNy�&�z�\t�����2����}6���u���Fe'Apq�k�<���y����4WW �E����?|[4	��~��[�Ĥ�.k�vT�$�'��/����+V���Vy�:��Pqb���N)��6ε��o7��=����$L~�L�ARBE*�Tf�]C��sYi�"��l�B6|��ka��"�X�K�j��d9)��C���G^��j8��ќΟ�}4W���s�ȭ\��X�����4��@b��*Δ��	lX��c�ŁyG�',��q���J�zk݁擏� �f5z��]M7��U��%���& Et	�L����)KĲC${��k���iG/u��&�X��c���ӎ�S/|�4�6�? X��$�'F�iϞ���2�=5?5�`�t�1IFP�5��Y�p��$�u����q`�ʉ-�(�۬y�i����l�_�T�_A-3�)_��%��m+x�n�9�j>�E"���y�\��^Jm�!�GA
�!���b�����c6��!�^6��>�N{��Ҕ�{Uv��i'�4/2Bb��Zh�"De��"5��f4�O�sy����Ĵ�_�b̙�&��L�eIZa/�q����fЧϱP��d^�h;.��n��q�/i���M�N�����gG��	�&��R��|���Iq_�_4��_@����	:�Kܕ3��p ���ZCCCenn&��tk����]�,]m���^.�#����"-��ƞ]��]Z���C�4	���Ҋ�Hf��"T��J�%��e]��x�����Q��<���D՜0R\^X��nx����ek(��Z���S�"���(�I���zjz&HN�RuB
�93,Tڴ4��5�\ܜ��M,��
ڼ ��������ˋ��{���v~��Gc�g�Q"M����&n�����=�.U�k[��;\pm��NJoE�#˕YD.�gZ+� D`+���c>�!�Q߮�Le�z��(���"�5��ۚ�Hr}s�YzW��`������Š'K<�e�݆�g����z\��u�$L�R>���������0@C�����S���L�����%}���!��`�ͨ]�����/pL��p���>UL����M^���PJ9:h1����z��8[֕�5=t�SN1��`�w�L��u����:��GPNLU���S�U�сS�Ω�>����"�A���#w�o�4��Y��v�x���SL噘@�[3���EO�Z^��D�A�>�{֘��Q�]���D����Wo���ld�cM�&#
:U+R'�M}_�^տj�:m���f8_6�LQ@��`G�+�a����ƽ�
}�u3iВ�v��h3J+{�E9�L���{�����zSʷT�r�h��>G�ίΚs[��g,3N8+�r^����[%� �h�֜�=�`,g�;��X~5ɐrg�.���I������fk��6y���Ga_�YMz�L���b_n����0˭k�p4`��Bk��y�	df�&���$�0Z�U�F1h1O�-���~d�^ʛ�H&�����"qF�wA�p�~������#�E�X^�䎩<ϗ,ܒ����b���%�\��l7�����J�o%�Ap���>*��<�i�H�"���Q�;�t%�ΰ��ta�,�\T3?#Z��p1.q����!Mn���gJG�^���o'ʔSS��Nn�#�����>U�<�"��Ebq�l�[�ɼ"��xF��������_�ʬ�=��j�����o�o�x�jQ,���|��n�&��5�A�J"��QB�����í	�QG�Y;��y�����	���m8՟#ݰm��>P�;��C�3�/�VNJ���C��)��!�
����&J{��S]̰�R�𹺰��y����7o�`q���r�Td���ڳ��U�9�ln~����Oh�o�+�>�qF���򓻡sM�����������n~�]^a�K_e�E�f�3�U�֐[Җ�Mm�;d���N�nY�ޒM��m ����Ȗ����]�K�L����m>�\3�;}�i6��s�%�&���ݣ��R��'��?",I4���u�7���9��x凉�k���ק�[$�I��Ǐ���_?�7p���Z��(��x�V����D폙���gi������S�"] ��x�J�1PD=�.��g����R��E�[3%������ t��컛N�����~?�o�/~��_?��Fǀ�KRf�53C��|���>j�c��T ������ܯZb�u������~���ܯ�X�
�~��x��[^�*��|(�����J~�yX��7�Z�&?c�o:���˴O�2��tR7�Y���~�7��ٽ����;�������/Σ2K�5c��D�<�}�s��⮙V������l��Y��*V�����f���\�x����J	�(����*'��X�����L��7V�����t���)�{�$G)Q��0��89��?�?����I���^�5+1�"!��T�������E	%{�䔔��Ay��f��{ފhX�\��B���vD��-�EH�̉�ͨe��ɓ'fP{�&ȳ"�m���cyeq,��_kմ���,/l;�r�d���@�i�]��_�ۿ�R:9 0e�N������@���Kb��,���Θ���x����n����0��[�D���*W����g=�b�<����E��%�S�ԭHN�DmN����M�
��\��y������-�&�&&��.~#�cѺ�w�[|yr։�5f`�޿��G �^�����[�,(Q%Ytf������;6Z�;d�����c2d�.�"b���8$~P7H�㨟,U�L�RۛJ�ط�P�^�
�|��23���Sَ���X�1��l�O�_'��~C5����|��S�`N���{�k�	�1��ٽ�J d��ꃧrW�|��'��!�7$����Gϟ�r�O����~�w���`c�t�F��7$���Wۼذ󷩢���8@Sq?)���� ����%~��Hl?�����4�16p�I��(j����G@,��^�:�g%�&M�E��*��\5���[��@��O�1���6���e��_��,E��g�9?C�S.h�5]j}x�kS#����FlX�	j� Q�r�A�S�9�E��\"ETjb��� ���G@8'� �����߅���z�ӣK-�/}�l����>ck��S���~<V�Y�'�g'�YZ�%�&_۹oiN5}NX���k�AUb���yO�����"R"�o��x��
?�A�Qi&�7�v��B��P�NW�+ Gg-�A��t�\��/�Y2��ߢ�O��7�o2�:�Z$����v@>��&����#2����X��f�iP��~)߮q�!���f�g��Z�ϖ2bsnDu 
V@o49��=~�6AΗ���M���%��%hRɢ�^?��g�>K��������#��~2��r�r�$��`���O��#Ӈ;(u�v��ϙ/�T�a��0��eO%� ��~�u!	)�F~��v�?�,CU�\ٴ�)x�+e@sQ�jV��\/�3���w�6u)�4T�MQ"��n�!�E*���nu����/��r�������$��[�O��SMs�V���΅����W������5�]�����߮��X��^"�s&�z������%�s�~SA<$Qъ��!���ws��֣U�X��E���	T������qRd�Sh����D~+�b�#rJ��`�ON���M9��/���U��2[�J�*��#����`3���KS��^=�z�`G�c͹?�K�F��*����G���,:�k>��jT���u��o1`���B�4jC�����a=�Aq�_�R[��h�j矕>�%���?��ׁa]i���&�QM��g�?�������&U���-M�סJH1�3Ԉ�C�*��v]�ɞ�>�V�Tx�@a��;{�4�����t��"�ۂm1_f����}��r?�t߰�;�S�k�[~����!G�����됈m�
݃��a3p='.^�Ge��Ak��37��Up6�m��e�h$Y \%S�]]��_��N���ӫN��䛟�TQ�C�+25S��k �����i��y� 29nG���a���q�[�xfG�Ca���:��L���s���S�����Bkߪ�!j0�G&@H=�UuC�F�mU;6w!��}�Ơ���6��eh.%8�Yҩ�N����@8�~�Yv�ʝbה�8���d�?b{_am{}���./V�*���̀�\�	����^�`[�$�a/�m�7�Ԭ�$�nu��M6f���� [/X�7����^Q���l�,�9χ�54�T��		�b7��jst���ߠ��v��UiH��>[�ӻ�TH�l�&C<7Z7`oN�Q�5"��a��T����*�|Ux#H���A_�yq�J�ҏ�Q!�9!��4��TL0LK[�P��^���9�!�L��-�-3-��oDI��ɭ�*�yz� ���9��ym���"��ʳ��LC�i����۩T��V�����D!���(n���\�">�ݰ
���r)|�HU݈[c1wG����=7T�Bp��L�>�Y�u��|Cm�=���Ɏ籍 x�T��m��U��9[7�dNR͊���z��6G����G�Π����8��ʮ�q�+����9���Kᅬ�U*%O�9����(�/|��j'鎰ۼ,�?�X�8յ 0�1���8�����65эΖ5<�:g�C�U*w��ٙLv(��;�nFR/hoJ&<*�kˢ۟v��#�:�;�T�VC�J�wod�)�U�L��b�����&ӛ6�	�<͎}~����^XH	��N���"P	b��,"��	�%�l'���Q��W�T�6ϜJ%�FY��
�m���C��#���왭ϔ����ْ�&~m��J�M����k���s�r���ֽGyZ��S?��@��MZ��v6ƶV�����̇�r<P���K~T*�����H�%?³���W��ÕXSe�n�ى�To���i�ա^��M*�[!�.�UPh[L�~�����u�==�Y*x�o0�dK@9I�xvU1y��u�+���(�B��CD�8@g�|N�j���ry9E��
��J�f�� �S����pTf�{Xо0�~e#�F��j�p�;}�*�ڴ3�"�((~�=�^�E���nfӭ��<���W�����Z�h�I=?D����GP�ٜ)A\�TCP-��}/fU���^�}����ԯ�l�YR�R�����j>��9��cu��_P�r�m�aKM#w[�SQ�MU�
#q�aG�� }7�H��֕d(��%�OTs�}��|�S�!j�q#���!O�1�O=O�2N��8ؒ���������nW�m*q/�l<K#��-�6o9J��-�9y��o����j����âm1Kl���Ïs��GWx����+��\�J_�9U�o
���S��3d5�\��g/�d��|�{)��OaQm���h�F'ء�	�4k���W��4S+��x�q���K�ue� �p& �����k�8����R���J�8y���k#_�Q�ʏ�����t��bX���=Sˊ�DwuD���y-��(��U�i�5h�c��i���3��ɯC0�\D��漂;���8M�U�u��˺��q𡾛�n�Ț��21�jh~l�a��-.�� �����P��M䍞G���^>۶
�n�b�g0d��ݚ7���ۗ�Йpd�k?�Dq�����Jl��G�d��6�L&V�#X,��8�!�f�O����xx-�`1�������^��f`oto��L|�7ՉY�K΋�Q�h�{���� X�U��T����Oal�{���
�r�2U�B9:;�����?HC��v��<�'�
m7��`s��f)ܖWY��YM�ԅ1y)��I�ؤ�e�y��X��YE7r3��F�W{��6����S\Cs*�9K)y�g��-ж�R�G���6��V���v�V���2/ Lg���i�������C	fp�P�:�Ϣ �u�Y�����=�º����8�f�ݰ��nK�P��#���Mo��� &>8{����K4�$)ޓ$��l�Ց�f�uo<KR��`kV�I��@�g��%&���r	z[FI�]).�l��)DX��U����u[�a�5Mǚ�e�����|JJ�Kq��ǹ�y9��J�������Hِ� ���q��e�y�O4��	i2�O��f"h�q#�Y�c��垩&G��������§M�X�E��,�GG�F�z盗ℴj&������:ѻ�b|���MG��^����`Q���N/D�U̧��hA��X��1[�ٳd��fs�G�Xf@o1g	��.p�v{F49-�2���W�1�kS �'hZ٥��p���w�����|!@�rT�'`���x�^.]�U��K�9 KI��{�θ�Y[�"\FA��
wv���f�
\,ٍ�%�a���V��T�4h�"7��^P��bt\n�w�z���n�q����,2YV�YRm������N-����gq�n��7�E/�i�euC�.�I	&s��f�Ω���/��Arv�>�R���1XD���5� D]ַl�^��.�1��X^ ���L��8�� �4����V�0���Aakn�p�|��Y��5���M��Mh+0 p9��=�;��|�K1��<[�[j�Qx/)�:k�	(�#R���M�{Ogd�! ʑ�
���0�������F��x_z���J���~�Û`/}iV�H�o>/�qHQ�����zy��y�V�'c�i�	�9��Q���@A�&bf��ԫ���j��=J�_6�~���FD~v?2�38^M�K�E�W	:2���J��^i�`�jd�M�`4�	~'2��PZ�Ո��L�`�$��f�!��Үԭ0���@�4�������v����m|RS*��'K�l5R�`���X_��"��SC����`mN/QS�ÊYp~����s�;��_V w��pR2B�h�l�'O��4�'Z7)�7?_�*&��Yʀ#o~�(#y*�Z�/q���7�_8��z�T��Z��y-'�[��M����w�j}󲝝N�D�G]%}�ed�L6J���G^+��x^G�� �n��Ps�^�I���K����u�_N�V�g'�1��������2g9z��p�y����V�H�F<��&>�۹Fo�.��B��F��B[�{�Hh ��Ć	Т����*$��=�Td0Ov͋���Ɔݑ��fM�\�$�X��#Z�3�}���ߢ�
$��6<�}s���	�Q��MP�V~��ޣ�e�:�,�� ���=Z��3eՄ��!u��1=ԫ��/�9U��H��ѣ>��}v��^/�S,�j�`.RB?~)���l�\�9������d��v�.'n��9�h��9ϙ7KΖ�.�[&A��]���B�>�M�l�$H���(�6�s�����`M���)�Ըr��D	���p����� M=��5��,S���Ț��5���^������?�, �]i:����}�~_{����m�w}�g���&�@���ݹ[Se7֠I](�����N_1|�1;��xo�h�ww)׮ݰ��Q8�f帡P���Y��X2v����9q	��|r�!M�2�n��c�fr���vom��*��a8!C:�@
�t5���nI�#ilK�p7�D[���J��d,�N��xW��JJ}4p_�%X�lU:c�lm��٫'���}�jS�bTA��G��'�.琱�_��"�1돣-�@�$���\���V�o �e��x�l���i���M�)����u;p�������2D�MRid�Ch�>��+�jS�s�������M\rFĩ6=<����_ʴ4�E�m�[i<�G�ﮱ��������@�ȢtP�'�x����)�F��.%�)���)-��X �(p�9'/�!����=JEF"o�ZN���e8��؎_I����1Z�p�5��l�w�G���;�
^+{e���D�%W�7��y�����}s�-�cd&p�]�X5Xwa��Ŝy���(l�dWGKV�h����
�W�C�-����k���"�Z
#6�w�'���M�����d���vF�@�3��&E�p�'3+�B(�ϼm�hj������ 9��S_�0�@����h[\�,�t	P�Z�=_�?ݕ!����l6!)m��43�;R)��n�|���� `,z<�X:!es�R-H@��r@Ē�J�KA���@K���G,�s�=C��EJ�N_@T��,W��Njʸ�$�D �j�lƢ>q����G��^��-�iGck�f��B�KB�\�����q�ZV��h*���wU���4�r�ĳT�蜨����	1r)U��Un0u�v���b��w��rEkՙ]�#Ng ��Y�p���"�a���Q������w��2�9qFU룵�z2��:�9��{�b��/ �^. j&g����@�U�f�m����8]�� ptDn�$��$�M���x��?iZ���z�F�o�ZC>���os�j�6>Kx��A�[ӿ�ʨZ�(���f��peд.ǭ�\B���^����[��-�R�~:ԋ�sW��#���~�~c��*��+n]��7u;�3�eOg�HV���z%��N6���37��0_uM�1�%��_E�m�e��CG}ESz���͉��}/?�D�Ci����Cԓ��ROt&�oӯo*���q�ɷ��h\�J���'Ăg
p��yBG}�y/�E#��h�4��%Ko
��IԹ�4)�����6I�R: Lي4��/
�x���MI��M�����@Y���iY[��C�t����?1C�Fa�@�'q�wT`���%hԋ�?08}&�f��@�#&"��L��ԅ�����v�uUp�bD.�Ҵ��iRh�&彔^�K�������	?�V3~im���3��q2R1����pGݷx���������,x'Q�=w��ׯ�t�:��K�w���s,�V�����/�T���ڣ��@�I�vqt�6���w�V�CO��&�8�l�����i��Y�f��Q���+������<��u��������`1��ڄ��a��V���]VU+���4\<�$��߅i����2�y�L�O�S_�����������(!�-%�P5�J�t�
���Hw�"1��� y����/♽�^��w�s�,[���K�l~��/�G�d*ŉ��c(����QFj}�)�.ǌ\�p\�;�+̾������߾!!/Ӽ�8���_e_��<"����\T���^���2Q���/�lV�\1)@��1�{JF�M��b��6���>ڼM�~~D��\�E��K����� ط����#�Ezr�}�D�M ���E�-�7u@�R�����Q�Ds�3��b0�Qe+~��CBqz=�g��������ʥq0D�?����^Bp�}��w�65�z��}9�r�6G�oF�8�U�oVկPf� ���@��`��� B��~"����[��B��k>�<���ܙ�,o;�U�w,�
|0})� C;�����8��q?��S��E�=GW�N��}��Q�,�(����/ҊW�!�d��g*~S�4_pX����(z���^f�ȧu�f'^f��K�Iw�.@����9�a���@��Z����Rw�0���lҩ'��y��W�V��O�r���8��g�4��M␅Ԉo�����q�����>ڛW�n�v�i��>J�l�K�=*$g[!���E��/l��-�����}_@�^=O�^
��OY�\8�!؂#�5�Jv²�II���gm��^�x�7���hx���ArS�*F���
�Ի^�Z�*\�R���ߏ�M�J[�0[*a����h:�K����P����*E)Mzλ	��*F2;�d�Iٜ��!��:>	��d��{��X1�3�B)���x����8�7-���wm=+b��a)�j��8)09��T(���>�z��J��3�N��dڄ��u�WpWp�WS�ٗe [���^9�H���R�d��핁������|�wo^��Վ�?������P�
���W֜^}xQ��D�$��.�4�۶n��Wݒ�V�
�>E?�ع��*��"F0�+L����FR�!:�T;GE]�Pf_}��rʍ{�cUG��%�13KF�i)<���n5n�	D��5�/`�ژ_�c���O�ʞ�v�>�ɸ���X�޷�yH53ݭ��+���zF%rª�e�Z"��Rے��<��K�����59����UG�ܸF�T��R��ڀ�נFA<��á'�*�t-j/`��X��_#|�l+u��BB/�%��B:���P�g�H������p�ꭁ��|ȝw�j&!�U�z����t����7��3?���_��M�/�c��e�.B�*���/ef�=�zV�q��t�WO{��կ�E8�3���M}���B������Z�}]Tei8f�v�vr��g�g�Q������	u­�G��H��F����Z(��C���K���X�v���.E��&�1v�;r&hk=D`�� �2��٨t�����7"2ƕ]�
�����_�����@`��j�c��6ZA�9D�p8-�Z�ܿ�ۖ-7��������7�k)�(����rX؈��u�H3O��]鈒cۤ����f���҃��>�"��%c1����=����k^GVA%�D�(3g8���g����7u(>��(?n?���Nv�I��Q*�]��EVfW�P Uq��䣌n����Ba�(������G.���qf�����czl�`��o��4��xyVj��D5�"ݲ�dU��v�x꾍�����'R�|�o1���O�`��!e���&A�p�!X�5F�[k��x9�5�qT��ɲ�s�ç+���c�*Ʈ�4�[�&�\f��}ȓ���x��j}�yZm���yAI���b�ۺE��c�������;X�}$�ڗ1b�`�ǽ8*>S4slc��� �Q�Z�[s�Sy��m��e����_{k��W5��ǩ���{�W�)4�H��O�ĳ!�޿����T�"���v ^yV��"#��3*N�炨w���`���G�ڥ�7,�mj%��bk �5!�gpM�&2^�H���0W�A�9;��N�\x@@�����Y2��F����Y"dJs=f���00~I��Y4_�/]��B(B��rQw�Rh��n 5���,�z�VA�uL=�GI/3i?J�r��i��؈b(�C0=��K��V�Y�w�n�V36G6�f�?�y/��~0R�W>�Q����o������q�"W�~�}H�� {L�ЕI$�#�O�!{[�n*��sWE��AFZ�]L\-m[~ɼ�$�<�l8�ݶ�A�?��גJϸdN�w?��.h(�z�NA�Ḟ"!�*)����u2C��I�M��WRv������''���@/U�!�#g,�A9qto���K��?��U��X�y|V?N�:��3 �H틠�RT[פ��D`�
����>��R�v�L�݋n{� 2]�*6�0�☤������R��jX��u�yk6B_x_�j���@���0�r��f|���m��,�"�ץc>Փ����4���5�p*9� dx~bWV�ýt���~��#m����!/��Ip;ҕ�2�X��B���!�	:�?*G���1XN	:�u|�B����%��+�/Yţ�\y�jaz�D;��K]$?��B��@�P���-����\�S��@^�&��}�m��V�� ��W�Ƌ/.�)�k����Jy��ӨQ���3���3���{��%,+ibRxq����"�$��`�C�0���Ļ�����ؙ�u�g�F��N�7$$ ��+Տ�)���@�M��{�j&,���ߏ
��U�:#_���I��ݔ�����;#��f3K��Qe�	4��7٥:wb�C�j"iu.n	�Tx_5[mV~<2d����~V�h��>��yf5��`�F�R�E����1�\Xf\u�*��~�B.���?�4!: S++8����$�"h���e���v��'^jc��}�MDD��� W���\o� ����3�yn��Ů���"/��Ik�y��#�c�J~Tp�����A��yN&��)i�S�Vy�"�؆F&g�/��2��'�.��`e����v�M1��(*S�9H2r�鱡7P]*[���O^ �nK_�6?���wd!���� ��^w�n�aa,V[i�zT�*�ȓL�����=P�Nh�]8��zICg��6����k��
��2��?�Z����)�{�^���V���7���Vn��� �o���+�h�pV��#�4^W�6ޱ���[�vl�W�����Jcr�KBy��2$�ͫ�Ɏ�t��硖Tt-��?fPT)�/:�d�f��G���;d�(�C������.��1�?����B�o��
o`C��%o-�	C��~W���?����֘명@9#!/ԧ,�yX��>�qgá�)B�F����T�<Im�~���E}�W��̼�tj�r����ܸ\��W�� _�K� ��x�_ˊ��Z�Z��C^{%�*�PC�d����C�庖/q� gΣDT 2k�ŏ�F4l;j|Q�)�-��Bz�#�bl�b�BJfhѧ�]��d�C�=~�vV�/F���e��РJ�0��w��%�nשp{ditw�[o���K<�V�����r.�2ˎ���7�O��8 �fɃh͎�Ӻ�l�D���gfP
�Sª�q�ԉ��b�+�����y��Y���V<]f�<C��$@Wޝ@�J.3�`VU^wA�F_�o�=�R\�nm�'3h?��i��0�*�6�z�h	�B�ĉb)���pu���j�IK֊��������|*�����}�eJ���)9{\����FaR��:�lŵ�\��y�0*T�5-�˹�d��7��z��PX��zT��Jq��X�YExjX��p��Z�BB8F|��0!�Y��u�P?ּc4�����˔�q>��~Q�f��PfGX&.rz���I�ѥgd��^o�1l�60�v�u�]�%@��8Ye�q�3!s��ѽ�'V��!ś�>O������ℨ�רu�yT:@b߁�}�y��a���yq�=)��@�J*wHi� 8:7բCx �ӈDCډL�[�3�
'��`���m8�>I�A��phu�ricf��a����e�@�]]�]R���g������({cN		�o��`�P^�42�;8��wg��*�;�%��@/U�JcmI˕�h:)$�����'��D���4쎀%7W	�'ۘ��i�s2�T|L�I_��/�&Za����)�Oo�y�8q���Llm���v�3�.��G���Q[!w��m�3A>��K��%
L�w��d�
�$Ku�Qi_���p$?��S�;D1W�^�#-|DJ�%�`�B��F<�F�uQ.NZџol�r����Fx�ytJ��RAqG�-����_�z��4'�B9e���i���F#:`�smU'sb'�9��f(�L��uB�X!-	0\)��}Q}�����c�!M3']c��}���/Y�)�g�}Sƀ�-�&I�P�E\��l/B?�� �m�Dc��x~ڱ�Г1UO�F��j�C��n�	��a_^����62��Sݖ� *إ;L@����:�8�� ��~�� ����k|{7�W�D������{��e�# ����V`I�R�=�"��Њ�	)�R������X��6�98�M�̻��cbL��y���|T�gD�P���\x<8=��>�����|m_�m�V�9CQ8��[{���;�i��n�]o�g����d�l'O1�2@��ѣ\��C�b�&]�y�� Hք:����ۡ8��%F_7��<�*��嘘9��L�f�~M�L=6�[�	]YR���sZϴ�еG��ϒ��n�;������闷zE�[{h��t_�@T�J�D|�7�b2;Ȏ)�E*��3���������(��'�l.y��["m��(�s�Ehɶls�Y��F��En����+'�ԤN�6-�~WQ���G>���N���g���?��a8w^�#җZg�8�K�����%? F�E�� �5�ƿ�^v �5�������}�#hxL�W8/���_����\��A�հ�g쟉���ЭS��;��Lw��g}p �f�j4�]U��%���2�9zn	�-y�����T�iu<軩X�7�j�_�c�t,$9���!�:ϴ��.�����w�>�p��Ҥ��!��z����w*����H/[e��_�1r�O�=����	�Zsט/��Zio��~`�TƯ�//xxm?l5]U@����R���t���tv�<\rsq�ԏW+<�?��s�Ր?khk�Ԁ�]�;$^�k�o�i��r&���.��{��`g��ܜ���ɩB�Z����3�I���.�Y�USS70�8G�HO((*��I�`��@��6%����onK9�@�f���6Ӽ�_z�e�L+�}�w_�c� ��M�Y���G-���8iu6�$,�݌#
�������yH�9XV��c7�F(N!�.��*�����cj[~�AJ��av���Lp�@��΢��S��_	���Z�;�\�s�� �o�<<����ύ�\x�KaUQʕ�>���S�"-}�XRu�#���T�[Y�oe�ѯ�lj����u4?E�q,��J���ݫ���(��5��e�N�|S�D�C�qA�����1FE+�K���S��K󁩲ah1��a�-P���
�p�qi���n��8�v%=4��8C	���<&���;�%���������(�j�0O��Ȃ짿C�$�>6>�c�ck��W�����ј�r�
��zŹF#��Z�܃�X�߇�&t-�=��-�X]]�Ze5u"[Jr�C�8/����4�����'3!O �M�H�J��G���;p$� �ط+|*Nmc� ���v����a��J�/j8�x�+��QZ�B�,�U�y�w�ĖK66���A�{��f�=�����N�h0c�xh�[�5e�~z�E�s��'��-/�%����-+! �X��b���4`d�+$��6���-R8e4:��yT�8��lg���I
�Za>�[Q����<\^u_}&�����+V��ЍH}��b�O���'�y)����:�U2�. 폚7���/D��C�<7���%�J힆�����׭���/��Y�ؠ�He0������a�m�A�����ec�l1��(�p&(��Bhu��U��&y'��s�������W����فoܱ	i����I.Ff�������ж���Q��S#�l75�|Ҹ[�6�П����D���t��q��s)�%����q��=N�e��	�ˈ~b�����g?��|��}D�'�b�p��]�}'G*������J������#�Z��i4�DR$&��Y��7$K�*��^��Q k��O�.�.�N�14����E��}&q,q?C����X�M�C2ŅŊ���2g��G�<:�k)��e��c��u�Ψ=:��δ���� T���R`�X^���"�-�P�o�1� m�aE�2ĩ{,�@|�n��=iI�С�)�*!�P,L#z�!>ݵ:Z�����$�p��(����E �|���f��������Wf���[�G�h��!ר�t��>���,�̐Y�0谕�����'���qO��8�}�L�8�n`�W.�7�ѮWqj�g|pF���o�����]�w��	��C�i�`mb���ؗ~t v%s��qj��{�����%�b�����F���l4?^��������?i���l�uP��bt=T!��h_]S�2D�*!fP|J곓�N��֥bgӨ+Z:��}قQCE��H�M���%:��	��X}��RB��,���̿H�y=H�T�KR=�I`61������<n�L)O坶�ʗsK�Uʹ�!F0���<�E���٭�yD%FUݸ�%���g��"�m�kܱ#ژ��m�8�xr���|ݴ˩ݱ�W��r:}������@X+����&?K��4%��+��7��卵�i�Y))SP��7��&%sln�u�ߐ��B�X1�{i��Aѧ��;�$ҟ�Pc<�;�v�+�c���ܖy�-�=����P��{��]�m��a		����j�+��dX&,{�>�{���"
t�^�ݨPl���@΋Ƈ!(>�f�0ZDt,&o�� 7	)���&:���U�*UP�(c'Eg��l� �������B��l93��qs���I2{�� |��S�h��^��n6,����4z��l_�M恛h���E*�̯�Y���S����3&����gm�a��F�_�QKx2)��9���M~��s�޵��0�9�v\�~ �����5�P��L��fb#bz�M�D�\��8�l+��</u���'�_F�`�QLO;d��{{_���n�&=�W6� �3=u�����1�P��0؛��gJ>>�����iZ�#���
C�j� }�P�å�5NX�-�{S��܅�����*��Eo;k�d[q�Wju��%�)�n<����s�Ə��w��i��K�,������lbY��j�̄���N8�u5╳=�����{v���"�-Ba� �5�Q�����E��Gf~^p6��q�gr��5�e��G�
��~M��d�Rt(�F���Z��wϢ��2��؉�0�6y��s	��༌ez9������ѓ�#��ϒ�E��d<(��飢~��K��UQ<2
c!}���k�wJ���jEa��g��@Kd�����&:�Kt0?����tî�c�q�ؑٝ����r�3�k:��F2LN�}��K$\{zɬ�6�Ȏ�^����%D�ҫ�k9B�h�t���A3��������^OZ�(����)�I�u��ԗ]45;T`�܊��j�|pu�\�f�{�f�����L&x�����̧�1�'-�CR�vE�[t?����kD5z����]���x��pɢ�3]��a�K��ԟ���Q���Hl��X �v(�k��%C��ͳ�ɧu�ͱ�<�&Ȱ~��;�!�S�(��G��k�s�v�^G^�FԘ`a9G�Ɉ��{��~��������ؼ�݂�;��}yV�>�,Y�n�����"��cWw-�+��=J��WBs�ZP�~����w�mƐ[na2�%��ƻrU:��uĉ�l��;��X�(1��WOu�/�(�?���
q<M�RwꡂKOB%G;��m$���Ҙ�zW2��̞�<�U����
ӯ�z��Ϯ�F���]]E��~�K�p���v�+ir�=��\ֲ��J	�^�)�������.�g���`�[�} �H����3�$��.~=�*a�K��ũ��(���~�_N�U�t�e��#k�4���Dk���y~��w#
x�z���_���KD��1�ջ��6B.��]|��/F�7��~	����&��l��-6Ʋ.�A=�Kw=�?�d��'5��Qt��H3˻}3�֌T�KB)�R�����:o��Q�/P.@K4�ҠP������"�dž�B�b�>�bc���:���k�m���g�=U���	�{��x�� ���)����5ǥE_�����'����ҩ0	��`�g�e�2���|�D��'F��S�A��/��k5�����eF���䕓t��+���z#^�����;M��Ж}���+Wܲ��>��.ZtAu�&�����8Po�۴+�ϗ�ﰈ"�<|9���d�g邡�P*�M���t�oљGtQl��íۀ[S޼��<�CS	Λ����7�5�z�7' ��,_э��R��8ѡ���I���I��'�O��G����VPYV3 �I��֏�����c	�8���z��ؽL�02�Ё:�d�g����y��F��3�Ӹq�5��݇,ԯ����8w�!�i��y+��.�3熩����v.�V/����ie+���Y��r��p��輥��Q���~D~1s�T�qo
��=�����"�� 1;�	�}r�Y���1�ЩSp�$�L�PCcx�����T:eh�����} ==>1�rt�!�g��vs���Vr��["�0� ;�~R�D�~��.A��A����Ö�.��_1f��
�dk����S��������Z� �&')"�-�[���%O����=6zHݮǣ���i�
WԖ�����.���Ԋ���u��ðK2����E1��u~w�T
�f4���0۱�p�z�"�$�&��r;X�{�x��O�L�*��vc����n�\�cD�^�n���2�Gk�C�2�����2�q�M���y�{�ۧ&z���R��Ơ&N�fǨ�ے��U�	�_��;?�WiɅ|=��^����&�z\��W�����sx1̚�ϣW�	Q
�6�Kkǆ�ɬ�aͼ.��%�zcn��y*0�+��L�0m|�y�2�F�d��t����\�
�����&òg̷Gkv�\�>����Y�.ru��S&�Z)E�I"�Ts׀�J! ��{̣>��]1`>�l"�Ru�q��l���7ff����[��q������m2�VN����Z��u���$t���T����d@���a����zc������Q͕@���E`ћs~#���^�
=��4N&��/PI�S#������-ݑv����i����VM��y���".�`�C�w��V�ݠV�L�lܮ���Y����&�E�*g\�/nᄫٝ��LZ��j�΅k̟9f�NO��������\u�b�ZG^?�Z��gP�/˾H�ořH�����q�3kͫ-kv%�Ɠ��p��Y��l��k\R�kϣ��8�X\�K�;(}%����&W�x8pN�6���W�g�e��z&���Ԙod�6�@`U�2���0i_�wg�C�-+�}�lSwT��Z&J6hZ���$�Rҟ�z�c@>��uO����DR�-&J�l_������wZ$����.���v��7v�	�L����H�=�T�pi<}�����}
�(�ڼb'2
˂�*���0p*#aC�q���{#N��� �-���A@}eLL�w��%������H�����?�T���G���
a��o�ç'�2s�z�!�2s�z1�/C ��1�2��zsm<;����0	=-����w�h��y������0����`g�Q��1���)`���>5|�;�k�k�W�P���H�o�\h��6�S�&'����Ԃg����z4�z>1x8�Ш#)��1�bi��Vͺ���Wy��󓋵!+n_T��*z�_���Eq���i��$4�~{ywZy.ok�Gr�a|~<ѐ��;����`���F+����Wue렓�p1����mw��`�,���{����ݲ���KUR*ifӉ�޸�ḎO�P(��Q��R��-mVw���M�@	�C �:�@)4�<�`�'�A�RG�.���ۯ!_�����<�/Z�~�f8]!I6h�J!^b�'f㐾��9�Q��E�޼~�Qu!��)���s_}��o����Fw0%��<��Gw�����ޣ_6��n擱��[wnȇ��!�R>�g����V�42��i��Ρ�,��j�eD6��
���<����w`j���>*�ȍ�˷�C%���o/��� �z�G����pV�|f���ϖ�"YN߮�|��cd5϶W�cd�Z����%R�)��_L�;�ɩ��d0"W��Ӂ���
�p��uDW�+uY1N�E#� �j��u,p*~�nd˂�
�d�i����VْT�����K�Y�� B!��I��q�K���;�A+Z;hJ���!��>[
U�0��W�2�Ic�a�U
[�˳�0�0,%*�X	3N��]q�k4��p̃��H�����z�+�o��g��L�^���ra�=]֦��#kS����-��r���ǳN�����ty�l�K��o�7������@$({���r]{��vh�{�G�ŖG��j������An~�^	[����������w�䓄�I�U�8n��Nϩ0����^q`����&4���w��Z�i�&,i��"��)T��׆V�ʩq��1���0@0�[A�����o �59i0*��b��Yφ�JS�+j��<y��Z>�����C�TW���~�i�72+Q�E�E���$o���^_�oE<�¼>��Q�z�E+��>)��I��{%'�p��,�:k u�31=��������w�����`�A�'���~��Y�b�_}w܁��ס��[��a2�Y��vCk����N��J��m8G�6�D�5d5�~c�nODD�@�=����%�PX��a�=��V{z]_��j[���)����ww�0�N�����wd�M�P��zR�<�>ܻC��(F%�/�|	�v�ˇi+v���\ e?X7==M���d�Ո35��B 4����˛�b�/$D���=���ΪX(�J#�����i�K�������f�Rm��7�x�;{w���>_^a�(|5Wrz�z:�)p�&׾�G�1+��n_� �tD`/�x����WwkW?{���p���);�`�̾?M�-����[{��^XnҦ<��8����<��y�Se�nmya�W�k���揖%�z�y0l�����#�v���Ĩ����,bI���o��e�A��w����zo��4�]�S�����1Ѩ�Y���ʆ�U�Cj�o��	u��Mk����jh�P	̦����I�/$���T��cm9j�<���Y�o�c��i}�F3�Z#=���3KB�kS�|��En�gI��ф�b`Vs]�h�;����g�w�mN���(d%~�vƈ���Ⱥ�{gp��_�}#��0�^�����*t՜x� G�SM�!l�LGSBe�s�m�)��vZd�?>�=��(��1���p���X�:�F���o�����z=�]�L��"�N>�̗kӿ"���F(͡�� ��41�q�T�lS�`�,+�\��{^ ,q�n�����^#�0gĈ�?���>�e5����s�#o�����!�4E�{Np��N>"���x��\tr�Ŀ����`^�Вt�45���O�g߮�{�0>����x���'�ISY��?#��7AXc�����.��Nӯ��=����h���~y�d�i�o����Vy{�k?��GFa�����h���0|�3��c����W�3�ǳy<��&sS�`.�k���������VS��`�S�|��Ͽ��  C��]%�D����q%���!�wfzٕ�l��/���'C�,E���<�٣����NW���%�Ч���B8�R7Y�U��E�f%h/�ް���ǭe<X�-�6�8�D !��s����!�!�B��y,�����:��I�I�֌�����oӌ����/U%YXb�6@���,"0W"����~R࿉�Gb��4޽��a���b"n%�s��99����K&L%��mS�ݜD���B6]����v`m�l�Ɔ������п�nM"�c��oS;���y{�V�{���f����!��%�<�����|�H��x��`�����z�������[6ذ�D
y|Hz�����v��~
�u��If�=<��g��t�����/�r���x�Sx��4*W�4s�D}�L�����D��t깺�Ȓ�3��Fc�!���/��+�%~�D/�]�g�e������eRm;�x�#�:>J}s���>
�P�%@{��l�G����u��c�U[����� {���ɡ���nvkgo�N?��ɝ=���(�	3b�D�����)��u|��%#����h �I�6��Xo%Ո��9��X��"��p��?P%��G=��B��N.��u{�t�	��ew��a���v���p�g�E��g���@�S�I�#"���?t�-�a�|8���ƍ	UaXW6����1�d|?����_{�?�:Ѫ�C!�D���"�[X��A�G�n��Rg�h��_V��h�>��r��9b�>��j.}�y�EȊ"�Y��, ��G��ԟ�y��ki�o�-j�sM��?�&3o���"d����)�=]����Q9�:�y)�=��2��s�O��M���VeT+yI�AV0~+��f�l���)���F�z,s �f���)���B���{���fX���I�����-��8�<�t�u:��7i<�2������f�-�_��
�����N�����
[@t,~�o�Sبp���b(_!�V��L��"���9P�i�f������3+����ƻ��%�˪|��W[�����E���$�ULy��TV��%F���v��Ս���t��IS5/�s�Q/��8Q�����p&��[�͉�����I�6I��U�������8��[���^�E�@P��+N\{K��8AEE��"$8��V��6�l"�-W�qXe)M��p`A���6VOe��aH@|��륀�e�!�m���V�� ÁUE��/�
.my��R��k�ʒ�:{)�[a!y;#��,G(�Ys�.K
���̌�<A~;������X�ߵZ�_�0�:�ܐ���^�}�N�m.���P��:�:wg����gz�C\#J�A��5N�R_�z����`�A�B4�#��t��y�**����������^�Qj���j��[��GU��-�'s��a��������W����aNQDT��ih��>}I��PS���A�kf�W��>�p*H�k��b9���p>g\����^�����	��NOS�������-�C-���#�Z:����=4?v� ��5-���g��[�I�K��2;.}6��ov/~�]].���s�B�gפ^��k`�<�e%�;�
�O�w�>3}T5�;9�*���Iݸ$�J�zE��/�(�"�K�M�j�h���!?ajy���i9��ǓN�}�^��LV�5�a`J�*����b0VG��./����GD��I8zF��f�BwK�N��e���G��-�����@�?�rB4)����`r�{�#l&~|Q]E!W� �������'*P�}id���ON�h-��_y��U�C�~�Hʜ �z�?�A���R�����U#���H�g���_f�O���۞@��NJ��u9qޥx�#z�ަM�[Xl�r,��-�
QHp�NA��2u ��#����V���p5@k`?�A:���r��Ͼ5߫z�^h"����,�^�ȕ���o�F|K�"�n%�v�j��fr?�%��;�f���ϋ���<���]>����r&��b���>r��A�/h�-)�����/�g�@!vs��[��/�b����|&|$Ϋ����_�/����Q0�	o#�P�J�K�{{�E�8'��W�� p�e����Q�
P�2&s���U�z(���~�T���z<��/j���$;��A�Ba�$v�2�3f'[�`����g91�)�H_2P��r�nԳ`^a���E�3�鍴��&R:���{0����r��.1���,B������)E�T��XԵ�?&�Q�q�+g[�_�,��x�j�Aϕ���]5u�����+zDٿ�F� u�Z���w�+��@*+k�e���"���I���a���R��� @���c� {S�n�ͬ�\7�9�{z��L��+�j��L�;X�j%tl�����+�$�#v����9I�� 0�d>�r�\�ӣ��22�+v�I�9����`��AX�xo�����h~���_�nX5� m-�}#au{;�k��q���۩���Ef��n��ٝ��_0�()�ޏ�c���6g?z��r������CfT6�� �z��px�5���}�. �1������� I�B��Z����M�`1�Ƀ^����Й���;g�:���E�9]@I7o5)ɺ�ɸ��N�N2�[o*?�
�s��"~����>z�k��Co���.�qP���'�P]<�%�����̻�u�7�۾¡�ޔ:�g��**����5%u��z�f�MK�r���n�##�sPE ������Z��0��ٙ����l�v{x��p~5����E��"�qҡ���B��^ ��5q�DE��$�F=�tX6�G��@FI+5�E �|�t��{��M�!�1}�^ҽ��2~I�����I�M��J�5�M���@D'�e�����
Ӗ�Y1��G�+3�b�L��Q���_������`��U�� �n�`��̀��$
�^HB_ ����ź(���l�}94���t�ꆠ�Ӵ:�@��k���I��'R�ypiY��U���א�Y ��}΂�\ikI�0���T8��O��U��!޻)w<����c�d��D�h�[{�Ts�|e/c�M��chy���pB���\H���*0��
����L�
$�ܓXy����\M-1���z���qRu[s�-��
޶�Ep�E3x�+�=h��ԏ�vG�x��ȶ��%�67�F/9q\��N��������*+k�:�t�Tଔ	(%��� ~R%�3ݡ�9�����?L��
rЅ��{��'g�ˎ�aR-���'�R�r��y��A�^��؊˔^��Y�JOȕ�?:(jS��˺��،�*���	s[V3�pP~�$�!�~ 6 l_����m3�^�<a���._�I�_�w�Pb�s:~��;S?Us���<n�Ư�{�UmcoV�Ol�vQt�Z�՗�.��-Ep!�XR_��\5�G�_�b�n�=~�����~���T)D�l1'q>$������s�C%�3��"��q����+p�������!أ)�O�P�cSf�>9��Fu����	�Lduz��{��>(��
���~J��Jϩ��TDi(Ց�eBfZu`��ح�Z��3���X4l߾w<��{�쌋y�y`Y�[�j�K�x>3�A����<���k��9�.d
�0���pOH'�����Ĕ��­�NdjT�����<�5=~2��Rne���-%���q)p�e�eQvW�������P����i&��z��ۏ����Bg�F��M{g�C~��y)�6�ӻ^�S�x��֖�;�Ǉ�"��'t�e�LA@=�Q'���t��پ�.ު������)�#ck�����MA�"��������٣_�/�a�U�ta�k-YB>_�ϵ��
p?�<6ms�q���o�\��br��a���1�A=h㈟�V���zy�\�S���#i�ř�A6�A�t�*?֓*�))�ew7���W�n�z�1����:f�>%��n��)W��]"q�a��Z��Ǽ܀��ŗ2��&��f��_�*Y�+�~7�qr��_]�WUS�m�Ob伈��m�]���� Q��<!���EWr���e�j�
�Ii�x�d�	R�d�TU���Q�̯D�/��j��Q5�����4�K���oR��y/��XR!{�cNK�wa�`�x�<C2��^W���+ꢅ��?���ŝ���?�Um��&��]tP��,�_�d�w��E�����Cq_�ƿC$X-')�8wꢺ[�v-=�-�����^e�Y�;:�G�tm ����~�9 ���/f��O@�;pXփ�)�\����_�ޗ�8]p��5��c0�ح�����66mf f�s���.Ms�q:�eݢ�G:�٫0�29������>y�G$6��	Phӥ4�P��x���U?�����./��Fη`�Z*��"�v_u������hh×ƅ�	@��·uZ�� ��`���M��[����h�~�����:BYz�����w@�-����
<�8�?]C�91f'�������/BO� ���ǈ�S��"̶�W����83P��ϯ�����ti.Ԕ��-	�D��n�r䩣Ɛ�Nv�g=�v����;HZ��3�09�������-q:����\K=��P�r������w��r�~�0����z�P�5��f{)��%{�[D�C=�^�|����j[��W�՛>��}�<����
��_�D�6o'����f����a�=��꺵�(6E@)�E�* �����HWZ��{�.�&-(H�^BQJ�MzhB�B(	-��p?�9�����c�{
{�5ۺ�5�^+I�p.��6�A����p�r_}KH�tz������_���ƿG�t�ɽ$Q6ġ����J��i����}��C�o¦���/��J˧T�+��doD�1���u�0���&�ܙF��܊�\{^�F����o��+^.Z�|dT��_���>��n0o�}^)k=��0�T�b�@sU�;�:�a��j��t㠃����G�'S���Mt��_�&��F�S��%K��.�J�L��w�eP�֭=5qrs�+�#�و�\�iv��� v������7h�w���٘1���;[��e0%M��b���Wg�5�ț�V�[d��Lϰw�<E�p�K;4��Kh�IO��}�M����u=Uz��xlS�����SS
�F|̶"���S��9+w�v�zؐ�^-�F0!�O�����$q8���)b_�N�1�M��p�T���ܯ�H���H�s ��K�fT!�F6�?;�N�Z�˘Өf��p�;x�E=\k9hE�n��2c����K���q����RbT���[Ʃ��Bx�X�ѻo.".YF�X�@���;k�_O�D�l���1}NhI�+�O�RX�+/l�2���)+�o8o9_�#��%VT��P�c�AMK�%cg����7N;�~��j�u�8�}�b�-����ӑlr������7�ނ��qf �F�ơ�tЦ�RT�MG׿��K��̻K<x
������;��{+���������v��K������ed����2h�5�)?�'LdF1�Y���p�jt��L+�EU}� �p���[+xdWF�&|޶=���)$��}w�W֔%Q��=g�)��fk�Q�eE-�t�C�Z�m�#�H���� ���e{���!E�q�˕�b:����Q�47_]�{u×��9�Y��q{�&�k���i�	��� �P�*/�(�qz�y�\2�/i�G=�̧5UIo�n�<;w9Bc���պ��~K{Gg3�t&�A`*�Q���-����.=�Da�l�*_Ba���Ժuv'aӏ��3�g��xrL��W�׆򱍗��z� ���Oc���k�R;s���ڱ�߸���(���n���)����,=K(�r�<�mG
i��.uu��ġ$3k���*~�ћ�?S����Og|u��ה��4&7�G������)��� `w�m�^Q�t�i9��O�ʭø����W� ��1ty�2�Lhp"������/u3}L.+�X݋W�׈��w���2�V>M���� ���1��c�f����R\%�g��+�T���Ok�!������H�D�ޗ@N(�z)M}�"�NxŤ��-�Z@d��\�짮�	��ƭrKA���0$v��1ٮ�~[}&ƮC9�եfƎ+��>�n��M�S�_�Q�y�e�� �D���{L2��ߔ�%܊��#��B��k;�O�@ ��R�s{�3ks�f�f�9�⨲A�WN7��꼢�����o�n i��	Ix�����R�Ӿ��Sn))���TC$?���e�H�'��BI��#�GC�v��JU�����m"�����ة��ML����1j�V��#��̌�A��ЛrF��Q�]?T�%��}f�O^:+}���
zҎN��B5�m>sT���c��>´��s�Ce�	�h��4���ttjaog��?�=�5g��mC;S�V��3��Z����f.bh�����c���EZ��3wb�
BrB�a������rM����P� �=�KU��[��9yA=�rSW�Wld�󥈱�w�`3-c�l z�Z
��,�)E��r7e�`fko���w�&wE�ĉ�3=������{� N(�K�kW����/Lݍ���ּ��6Y����2��B�%�`���(OI��'�"����B�{��}tf]m�E�u��2@�����:���~��<�>���=��������[�a�	��z
���-�8����8��Ϟ��}�.��w���Ȁ�h�4��;C�L��Hf�9U��ʈ�<a�ײރ����Hެ0"�EVA��!�9��e�K\.���w��}��7;�V#ʺ��ռX�X��8�fXt~�Bh�sI�Ȱ�pBM�6K����A7� �H c�T���`�K�Q�'!��ŃZ�l���˟��-5wDe��C/��0��@�+L_�2�MtQ��-h P�����8�~S���/�{���Z�qGG[ͥm|\�t��P���o�b횣 ٵ*���	l����p��O�4����e����=`pZ��ǈ���?��@��@���K��}	����vG���e�#���>��M��C�K�q �
e��hURm A4�ݶ������(Z�k�N��:�;��7�ΈT�"�:����>m��|��ɑ���iG�=tw�&0=��)u���ڡ�O���1Z�$B����*��o���g`a��������5*����b�:��*�)�6�dB�Z�b��xb�����d@O7�X��on4�&:hS�J�d�e^y�O�w��$MGR��Ľ����a(p[�	]��J`S,��0�ֺ�Fzb��k�{�?翌�p!l�����8��2%���{�Ivz;�c��]��f8��(O�o�͝�8X��GO�`��'�l��8�h���i��/��r�
�`?^����'n�%A���g@n�G�

~�uE����x�(T�U���a
��顯��1�����ik�\���H�F������.�ca�~~����^��2>�8�B��M��������H`�ͫ^�ǵ�T��1 ��t�
S��:y�t|gh҂�*�R��#>4����@��nT ���yG5e{�ބ��;	Є���:ީ��}�T��!����4o?�0W��8�ɣ�Ҏ/����j��J;���6��6�~W0�o��,+�<P�1o���o�Senm,TF:N-p��&�rTu�_�!�}�#`�e��1������ՃF�Bę�q�a���m�x��'�~���o�7¤,M�"�1��b���*x�A�_�W�x��Dp6l;��x�>���F����z�F�������Tb���H㒻�s�'&Y<���<܎@<��ÿ�q���������{,���	]�ݸ�!u�[����5��2n�rb���	�啪>�v�+?�,�ڤ14i$� �"���)���"��!�?�^i�����S�=��o��vd_eٴ�f����`���4!ce��4;?�,�+��[�B̘~��OX/xΕZ�3�'#%�x� 6��	\5�ca1[Y&�gy)����<�OG��qj,����
V�~��)�O�kIwN k`�xOrJZ���bǥ���aNj�3�F�-���'��Ip�뼮_�*����_5�D�
�0��'�_�e��c`Ą��'���v��(@������\�+�kD�d�����t"*�c�F>o�t'���u���yE�s��1XN~I�����u�Tɓj$
_f҆��vD���	N]�b��^^�xUD�*J�߿�y��������L� �>1���4��}a��C�����)���S��2�S�J��/'K%9+P�31��|�>�q0�(�<U����Ǡn��FeZ!����T�ʴ ^dx�ֳ+�jӅ`��a2Гn:��Lۢ�g1���޻�������w�H:���h�4J�}���lk����Rx�R�����Z����কS��|w	ʿ�Ό��~���1*ܾj"�.3���*�d~ (T��gKrlG�cr�5�����
٠��l��
b���ܲ;�P���B���E�/B�&,�{�(�4�V�u66�^�{(��]�>�Y��R���ƿƿ��F�{dw
��#�E@� u �%e�WO���9�p�0�u�L.;�i 8˼y	� �g��! ���80��@e�"��x�P�6��e&ju��o���^�<tt��c��71�*c���>C+r�l�ݹ��X@��0����ډS�ZB�F�`^���;@�<݀x�-8zn���R�����̳�!���$��7���o���<��X����
?S\7{Q�}�uO�pv��očtK���ȡ��c��򙟟��tR(F7�/�/��'$ᑯ��h�ς�s[K�
a���� &�U��U�{MO�=>���
#;�;�v����1���D�£ ���5j��Kn�t�}`(P񷪲���:���GV� K+7��cю�XxhsZ�f�5C�}K�3 �nd���A���v�Gb{{�B�Y�[5-�g�aY��Xg�%t^v� �(�1��tթ(��G��ãe:n�U&���!<(�{��w��Ռ
jD��Ĕ?����/��'��O*�7�
�_D���7Ӓ��`�:��VzuV��,�ʷ�����ˣ����K�������\�rE;+��a� ��#��9߃`��~��2�f���dP��5�&��I��F���~��A�+.�U�Q�y��B%����F��|���yT���^�5vM�Խ�NA����M��Q՝���"�|2�e�Ԕ�&5)�a�ëj�4�%��2�������I���M򔃭ߟ=���i�U`iE�c\
JxIЋKUF�UՋ�<�-+=K���O� ��Aa���މ�������I(������j��k'�
]�Ry���VQfyt]lLf��Y�H�e�J(�xJ��RtY3j��:�>�,�'p������DNڴL�}�mi):��`�>įY睸)����:�Q.���}4^n��7��Y���;5 �&�(U ,"7[1]������sޱg�ZnGj�n�gE�-E+e#ώ���$K9<��0��������x��[�Ϫ��S]`!"Ȼ�������H�&� I=11��!�gfg����"4�ڰ\N��aR&p�8���d1�L�q�8�1O������'T�c4GS�Xn���F!��H�W�s)���m%��R��	���4Ϋ�$ى^�s���_oPՉ.�poA�&�fղg�1��Nj�Hy.�F*�͛�z�8��q��R�H��M�s6�"9���|���!z}'���N̚L$VSW�b�6�?iG�Zn���e&�M�*���j�:��01�e��pVدM���*��#��K�3� �d�qE���=�CV�)WjU������Xc[����֒R��>�fi�)
�OȦN1��Q}3Ve�޺g����RÈCc�U�h�D/���ܘ��r�S��uz��h��f�����e�}���F�_}@A��F��p�s�%�����V��G�:���3���4��A��,�+1�L�_��H�sy��J���{>F�H ���) �����:<�ٜ�����+%+� B�h�O��:+y�@�$Y+g,**�*a���(OVA���f����nF�$��*,��(���[�^Qx�l�u�	���Z(o��C�}��%�o�	��Z�8 X�
�����s�ȓހ#X���e����}���{'���>�(7�w��ϗ$��.aV�3�]>��[`�rͿv�(��38�cy���` �۲m���k�M�q�ܾ�*�[[�-Ubf���\���Ϯ�+�`��mR~&2�y��K����7�B�K�E��,����g����9ڨ[��fő��c�S���;$Ȳ9�y�p<պ�q���r1������c��kVy��m+Ӯ��Q(af�YNt��7�	\���5;��AF��vϚ��d���a,�Y��T�Z=�����>|�}f����Gj	2�DF�m=P��iD��D�1�O���W��FYĤ^r�fQ�G.V'~�Ŷ���\x��<�)ѻ�P#.ɑ�u�-���^�a�sG<�vD޻p��~�T�é)�m^$a�߿�g�N�m�[��*hI䶂����6GD�}p&�P?�ޫ�h�����J��*#s�m����UE���m#��pf�e[��*�讀ڊBq1�	z+C�~���
��j�W�Ŏ���v�G��^�+3��ٯ��ʉɽ���F���!������I&��x֘4z=��Č��(�)�@�Os�;�����ӧ���:ڡ$���˝�4,f��suQ�g.<{h[	N
u��U��Pltn�شٶ����u��i�:���Șl�0�+��W��x@�9��7�{x}�z��]|)b_�Ք��63X��y:���0���R@��ٻ����])f��]�ŕ��5�W%,�e�M������>��{ՠ�ko����������Gתkl�������$�-�վ���7R�]IԺtYP�O)W�A�Y���e���ќ��D_�eaTa=�c���k��UVN�������梳�l��������l6_ u���y��s��w?V
�M]�L�{�$^k�.�� -�KD:��f�a�t��7�[{7��:�vEs��ɡI ��+�2�3ok�{�Wv�������Dp��n��&�Ȭo-��+�����+�V:G���C�BlYot ��EU���J%Q�`�Sc½����"+ܬK�����xc�ۮ0Ψ���#upf��]�0A�iM|�>`��-ԎC��5 �ލ	�SU���e����z�ʓ�@amj���`����z�=v�WZ����]ގ��Q�dB:uZ����#u2�t��6�$�������ͦ��(o��G���㥦��6��ZB�d�R�l1J�H^a��<z𫕼�õ���ؑ�r�LH߰��l�1a�S��k�%�����j�N��.x���b)�G���2�q?8:+�fa����{�����L)ˁ/�S��ܢ�f���΀;�2�y��ǖ��d�m�}Y�̣L�gcľ}��ꧠ��ƪl+筹Mܺ[���A�Gh(�#�*V�?Hx�<A��W����>�� �'h���go"�7�1?��$�4⒮E�ט��l|y3����iZ�x�ggƃ�^f#<&�>O���������U��ŌEV4%�?�ۮe`��0�@ f�坞+�Y�F���n]M���:��f�i������qo��;��5}yr�M_���zB�.m�����	��[Xܱ�
�w�+��hltƕғl��j\�.�_�u�N���#>4��ܺ��+�F�7��.�GD�o�m
4x��]UrvRn�ֱ'$䳬�i���6e�����k{��L@�����AIt�� 
��f��Mb=[�F�v�#��e����u_3
��R�/%e�LG����iz�woof�@�������Fz�6�%M�T@��E����j2���̲��ݬ��k�rl�S7��B�o�9����y�w_����xJ^��*�J�#�m���`q���;�Y�o�d��[����m��ߦ��o�$�z�'�I�h�B.TPL���T�e/ڽ�7��S��$_t1s5�Tńu��Xc�Z'�sS ?�T��e5�%}��?�Ў�j�&�jj�>���"�Z��H��&z��_�l<�&wg�`�n�n��wQV���@�,Oﲉw9��M�x ��O<��iQ����.c�[���o.}D8��uu��aK��ߎ�,}��u�7�Ƈ�H�:j��oom77��D����I�侮�E�t5lwI�KE�:���v9'�/�g{�7z����"�� pG&$5ƺ�h��C�<�H��Gpn$ �l���/��4� z��T�w�#a�aa@*��ܠ�~.��⓼)�d㿽{D)��m��mW5q���i��`嬞|O�/��<F�~7&��N8����24]� <(19����v�+�)/�.x���6�鵚��eIiY����igr�ߔ|���]hiE-��g��������|{�ր�c�"av���	��'g���R��T������d!k���l��>u��1��
�>Tj�I��s^�q�R揘_���U���n"V�D��49/�+1n�l1�1�0-�S*�;�2��4pһ�Gj�0a� �Ӆ6��oJ̙�m�i���V a۳�hs���
$u������1�?Ʀ�[7��	�)F`�ۀF���5/H�6��V������5b�W��.��?$'��*U��'lq�|���L}��!Q��ަ��|d�&z�����

fP5>��/� �6��C
/�����lm��ٵ�ÿQn�~/���b��f��l�Wk�l���}F��v�E�t�f�+m�xӘ�4^Xk�#��ҥ{\��:%�ݞ�Q
�G/Z�q��,Ք��א��́����ʕ�F1�5\�&��@v�A�Ҭ �_X���l���x}�p��[l5T�o���"��˶�������w������=x<  d�De㻟�Oa�c�E�I��bN/�5����.��%(9Lڎ�xP\��Y���1E���Ov	P�x��'	�]�i-�_��tk݀��L+V����M�W�U��}%gq�m��^ Zdsf&8���!��%O���fi�����,G�U�;��eeŎ�%�DL˺L��D����Y���0w'��a��据���&c��Ћ�%o퉾>�6~m@�Dl��e��q�Y�8S&�R��e��g�~���}�m�t�J��B�Ծ�+�]p����b�\�%2�N�dȭJ�Zl��>��EEhr#<�+��PuC�#Y�'��5����o��~�Բ2�����-�C,�ⷹ�˓����æ��7^��
i�L�����9;���$�9G9�m����e�x��՜����We~�.�����k�]2ΰ]k���AZ潐d������a$v�Ij�G����vT�k8/x�!|��%�ze=:�WZ8���d�Q���b�d�c�Z쪓�݈7��DS�����K+���3X\rZ9�, ��_�l�SjTR4P�q�>����*�;��	|�s�|�6����|(b��eAÚ�Z��X���Iq]��n�L_��:!W}d�(�����8z� f�k1^f?i�/��4�dSU�,��޾��$�y���n]1c�b���g,�+��L�D<ep绗҅����Ѐ�/
��̵Õ���{�;��V�@�%/���O�0A�NTG3P��+y�o��UJ�����9g�S���m}�K�.ۙ�BE�AO4��'tJ��⢲΍ q<�z �3W�Y�w��|�%K��x����ƫX���>�������=56���w]�����&� ������z|!9!���3`����S����nƒ��Z@5�g"�]����x��'X$�7�)r�+�2z�҇�\�L��b�R�����t�¾�5v����C�.�|��ĠA2	2t�_���;���y�����ϔ���<���@y��3�Dp)`l�|gA�=�%��Ldu|%l��=��z��g��]�)�'|/j&����,~�2�ɸ����K��]#���dk?d�؛����{wM���uq<`�w{�/�߬f�#�J��1�� �*\��W�� ���g��o�
Ͻ��~��V��B�X}������+m+�(˾��do�;�Dpp�8��3����R	_H�$���2*��Op��ppd��!j��c?��n^�&���1�����qV+��(9�U}��fO��RM�R3k��?��&�������HhT� �v����u�bx��C&e[�O�na S�T�X�W�+�s�2���������~Cz/�`���&'-��l�XH� Yk�*:	���*���nMڙ"�X�ό���ϕft1| S���;�#���%>0�i�?j��cRp�ላ��tD��@IH��h|OKc�n3�?�Ԣ�`���]��}����`����h^��8䫡@�K��@��w��z
,f���B��)�s���8� ��K��Q�=WK���@�Q�^Q$[}Po�K:9��j�b:��R;��*e+6���T!b63[J��v$�DN�̇{|��a�����pM�g�>�ހ��������������m�Xd�����r#}�䵮�X۪4_��Er2�^{�N�.j-H]���rK�5Ւ'���+yB�c/��r.e��@��U���U'�ؕ��$�^G����b��1:���/��f��2�OBLמ
s!#�5{�l1�Y�A?9��r�w04�n�{����䕛�u:��F3f�F#iC\!��>��@&j�>�_��;3̠���4�OGm)V��^F�8�fU���\ ʝ
\�aͽtHQS��j���w#�>�E�/�F�M���g�r����۱6�[*��6ĭn���]<3�Y0F��=�I�\˧/��L�������6L�EX=Y&�xFuə��E���ա*S���Y��[s蓇��\�x��'�plxH89����u�U�.�+�Z>�i���9%�2T	Ti��XqL8���׮ۣt0�f|���q�,���$%�I�H'y^+�u�F�z攡=!�i��Uhn��5��R=x��ij��',۹`P�� j�`��$'���Zıi~�!���������W�'��"���~�7{�i ��H�� (�{S���g)z��� ���Kv&br�v&��}�i(�H 	��zm#���?� ��������:�yX�rU�Ŗ��?2e.�@����������oHb͑�z�{���P��,�]V���J�`�8� I���6K ��N� c�U�L��Jw�1��uT�V���6�����T�ZZh�p�]!ynj�T:�~T2 ���Kg�R�-���"J����t?n(���2}n�@߳2��f��!
M��+�1<zXI���_�n����}�*���4q?�b�P���?l���ܴ2 ����0^�uW:ᥴS�`j�a�;֩@������)�է#�Z׮��P�/ݡP ��*T�"Y�H���wĆqA'%�O��}�*�f4�֋}�,9�˗��yz x��ּ�џ�������@r�c� �v�$�S(��gg?v�^�t{P�5>��[���m�RuQ��
o��h����ъ9�ߠ��ϪW}�j�M�!�{��4�GE�I-0�&���}\�S����D�#]��\����9�"u6$�Y���1.��_��
����k�X�V��Ki}�lV�� hQ�eE�W��T��V5��+Eqᮚ�?��>�J"���l�W�i?��3��4k;^��JI��Პ]�s��O���J�,wHb�t#���PB���
������t�&}7�
 9
����-����~�[V�P�ɰ�?@��k���g�AI{Ys���0­�V�H�=*֓���O�YC]s�ܯ�'7�+�"lN��
�� ����690#�[VmA����.Q	='ߢ�G������n�ck-�W	-z|<#4enP��_Ed��(�U���'O��8����t�w�{6E�2?�������O(�,b�_Jӯ
bâ�1g1��?�G� V��i_����G^�#?z������2��� Q��]���G�	�6}}i�u[���쀹��
���G:/���§Ji��vk�����;O��e���6Azs�D�Hd���'��jU�"��������)�ހ]���j�nA�9�wS����[*g@7�4�C����c��mW�#
�k@/��x�A��=jq� �c���YMQ�����\��%�#�(jj/���v�u�St�dLT)AG���dHf	��F/�,cE�3�Uܼ�|�9���k���jN[$��T�=u
�H��ob�s}DG� ��k������	8�a8�f�(:$"�x%V� "R���t� LT�E�p�2jJQ�o�{�	\��'���?Sej��Y��³���Q�aI�:]��>�.�>K.y`��hYeX�!I:����I�O�I���~j�ʳ���<<�}��l�i�k�.�OT�=/���.�j޴�1�__��!��|$�J$�����74t�G��]�b��ث>$�/Φi�͘b\�Dl�iJ/�CB�"a��,�]��Vf�M��X�4��a�t�~��]���{`8���)))�HpI��k�EئїU����a�Z�w��|��Q����C�B���)�xl��'"'$d��S�Y���~{��U�+=�m���Gs%7�,֛���*�|�;e%���Q��=����CII�Ii�O8:���hU�3�-[yކ��[�Z�����gU�߄�Jyמ��Lj$�uH `h��Xs<O(΍!�-F��Y�f��Gj��N�O%&�/���\���P@�E�iϻ�+�n.mZq.����s��T��~�	p�åါS�`M�_������!�ri��0��*���|����e��M�dY��i<�����,˘k��Ԯ���#����Z�8õkRs���c��u5�RR0����Aʴ�����E���M��V�����2_���h��֊�9�2�N�~�c�q��ب������Ӽ��*�B���z)��0�.�<��7��aRt�3J»ҝ�K��,���)𖀼��UM�d3��*(�nH@f��d,�l�2Lܽ};�%j�-���YEƟG=H�2��O�.�y�g���1�M��N&�:�ܐwaX26%¯N]%d��쪹�3�P�UK���'�7��T�&��o��<��_�Műfe;b��:'�7פ!Vo'l�T�MҶ��C>K��脲Ć~¯��Z3��F�-w( �)�|ܶ����Y,[������z����sy����Ƭ�f�����(����\A�p��0ۄ��V��j�^F*nL�����S=60�5�l��*�W0�|רj��">��oc]��6�4��]�=V�
�j_(�o�H���| Ux ��_���L����zm�X����޻��>�#���B��I�cke.]n����ڒ�(��4	��-l>V:u/&3����F�D��Z����5g���{�Xc-4���Q���4N�1��d
��\��ݬ._n�I�v��}d?&������K|\/[l�Z�|k�P_�����x�}�� [���Z�kO���1��j�V�s����=f说�-Ȥ�K����!�F�����	fУP{�,�\gv��m��E�JK竈o�K����D��ar����Ƿ�'9��o?cV���ap[�*����,�N*�y������OBZ�c��b�f�������h��\����gj�^�B�H
#x�k����K8���Z��`ɧ�ZW F �
y���e��>?R6z[���Wc���;@�]�dvB�X���)�B���~ҳ0�YY|>	~5B�Z�.߶���dˏL]� m�i���g��察OȬu�30z&���R����)����G�g7�g�ڒ��(���ۘ��M��~���F7U���L�.8�ߠAN�۞�Ǜ�+�WY�����]W���Z<oH���I�
��ia"jU����Ϟ��N�@0�ݸ�`���^��nNr�4v��".U<��>Dު�-W`��p�G�����9�5,_�'�A_��d���BOٽΨ+i �v۩ z�6�M�pg����b��@[�K�C��䖝�d�M�c�c�j^�:�����j���>vDO\)�����M"`�u���\��ѷ��U��bXlޥ쑃-T��e?�|�f-'^j1 dV�R�:�Éդ"A(��+"4)͂�����p�1z������B��W#�N{�P��;�'�dc �e���]F(,d✅�/���?�0���a�%�ڵ'd>N$��`��?���h� � �� �ϛ�63�mi��	��*�A�W!���
'�V����,��֮E�k�C�ig�a����4�U#ohڝw�f��B`I=M%cS~���-������K5�o���`��m�>�,�xL�?q�ߩ�b���	�c�L���	�8�O���It���������o���'4\��SB�I*J���
���JI�/a�ݔx�6�W�IVq�7h��3K���W�����U�� @[�&�t�U���PV��~<�6ꈘ�c��J���L�~��
�:.�ߔo�������g^e�Em�����}�B���>�|�	}>@A/�jȍOb�Z�3���[ҡiĽFg���GV^�!�ϱ�:��8���
������q<�����gY�?�Qo�<����j�7*��)�/���^�KWR�M���֠��&��i��/2_~�z�T�sI_����U����9�cM|u���*%fIx�]'��qol<;�����HbYL��c����9(�ZhRu\;ɳyy���*��%|�XC��FJ� k�_Y;��)�l᷀�S[��.C���#�� ����+}S���]?���ɪ�3�X�Q�uמ�`&�0���- x2r+�YƸ�	����I��=%c�˲���yb�'[o���v��$�*+M�Ae-T�C]�hњ2k.pf �b�c����V�r8:6a�ݱ�����~}7�����9�����qڸ������.;�s��v7�"nc�|W�m��m5f9����� a�����aR�ғ0���aoAM�D4-QF���1`9Iz��A9�h��*<5�~|_Xo�I��M�%�Sv�k?3�W��烏�y����	��냔��3���)�\m�� ���L!xq��JPWt8X��;�{��𾴃AL
%-�H�����.�G������>)�0*+���eߨ�;�.--�lB
/�m��V{@J��V
]��Ӄa��px�=���xLg�\�\��L���;b�dge�t�8P(�?3��%�dR:Z��M2Y՜/$I���֕aZ��$`� �lK���ۨR��Q����?�$^W�K��<j���e�E�/�&o'��w�@0���y���Z�!p=�^�T�x����������w6�[(�{Z�qp��ݷ�=,���ö�����\rSԱ�h����r7�,�y*3n�\��N�=���]�V�>�O��:\���YZf��<w��ɲ��f�� }{�Ԁ�Ns���γs���>�!��e�S� �E�Z-x��
nGk��Xv���s�^�:��y�I�t��Py��Ў�b���F�J+)aFB���裏�r�I�>��ٔPY��U��b#��b�_d9Q�����juu���k�]�o��e6V�b������X����O��\q��n
54"k�-�t�)_�U��q��@Mj=�k��(���2,1���k{��� �f�?�v�ɞ�~6G6ډ�.��k7<��E��,���p���yI�Q\uSC,�eZ��"�{��;mm����e"ߛ.��%|�c��I��0k�}?�o��|���j��Y�)T��a_z���l6�1z�C�������Ac���E'��XX���C$y��L��N ��;q,�qm~�݉�����t׉�	�L'��@֖��,�N3�{�~�(����y�N=��g	&5Ǜ�ŕ�N_�������w�N2L��~�9��OP�4�cG����k|��=�VDW1V�;�j�Ew���� ���
�
�O��]�@Eq���SN�$�;�'N^~����[������CJX�m�E���uw&��\�,c�g'�n�/�{6��3v���m��WVC�v���%�~�(�@������s���r��=�N�[[����=�ӕ�=��y���Nk�������rG֤�5G)Ij�)M>��CÏ�f�q��n�7���'p���P�x�\n��#��tڀ�����L׆��g���*<\Ɗ5Eb�=Z�p�v�J�s����z��a=�+��	A��NOX��Ȕz����c�2�o3�zf�Y�8�h����Ȳ��k�Ξ��]<��J9ڎ"���Tr��|�%�0���I�+�Q���?�8Z^��X|�ǟW RG:���&@�Cצ�M�Ҏ���5��*K�a����v�U���i�l�yc4��N!TF�Ҳ�v3���z<�v�G���3$��l� A$�81�)u~����~^�k�k!mǇ�k;葭��RUުA��Ѥ;�r%/���_a���X��g�3u�^Ѳ�{/ :z�(ޝx��{	N"�v����v�
�}��'NBU������5�{���<9r�K0����2ܕ����n56���D��H�`*q��y����!)��~�w;V� �K�.ci�HK�_����Vrޘ׽��R.8@=Yd�N��)�Y�����?<�UO%|��e�l�%`�w�T:�n�hI��f��4�p�Z�d���&���O�����:{y�8����1�{�������Ƴ��,Aۢ�*Q��5������u�����-FO#V��Y��o�|���V���H�,��^������)��[�\�m��E�Vv�gq/��%�ڬe���S��K��W4;���"��}�������<K.�8k�S��g�X765?��^*)�� J.����Ը��7d���|0l�Ơ�T��։[�I,�6ڷ�J�P�K5�������ק,v�g=W� ������j6~<iuQB��Eh�����x�Փz�78�s)�i�ٺ�j��5�ξw��8����n��]�{��������A��K���Pt���'���^R����u���;�����_D���D�"�(��'�,���:���/�����@�/��g���O�x����+6M7���	�%~c���0�,� -.��ȟ�p����)����ةb��Z]}>y���э��턊H�����5�Ȝ����u`�I�+b�u5���e��	��"��Z�Q܃EI7�����j����ߵo��m(�h��Mr"��Z��ᓅ�d�v@@]�;`Ƽ�2BN�U�c��P^A'F����E���Un9�E`���_/���MY;�����8�o儜�jG���~F�(S�,��.q.)s�c"��^�_�3I9��Fu��s��O Cרs�k3���n}R��鮺b�,>i��yM�㞘_����0>����}�		͹{i�v���np����9<v�LN�c�uC�i�t�ݖ�o�e�3���E�x#[{Ə��G1ՎYs�*e~.u�[> ����U�޽���Ja��J�&~
����K��	8�h��3`z��k���R·�E���#3��k7|����5VY��R߲�K�,�ю�"þ����np��?�L����/��H]8�g�t��S��H�^րK��e���9��,��Ŗ��ׯ��r��;��A��8�Zx5�������X��Z��jǒ��/�R�Z�d��k�2���f��˾����s�
.u�%y:�ynv-�W܅|�I.q�X[����\��j���An�ZXH��O�sfy<�wX��/CaIesAb"�1<Qf����h�갦��}Q�RQ:%JHI��@��5��K�D��a0PF7� ���Q��ޟ����K�:���>�y�ׅR�n�ǻ=�JJj��h�r�����d��4��!�+kh�ҧ㨩}�㤑pr��OE�E�����o6�J�' (^gY2(y�U;P��4�[uWM^K�l2':���Ŏ�-Wާ��ʶ�/'�EP�w�B��׽�8S����	Y++��������J���6̖h{&),�����0��_�?����z��-��	�:����6k�;�v���Ѳ*��j�cq�_�Z_�o��]-�Aށ#k{�i#=(ԓ' ��r��9��_+���8w=�0�FE�ΨJ=`��LW]1��᙭cP��]U{��%GLLK3̐�=5V��Z���
���H��<����SM��ޞG��๧O�?�����Դ�Lx�v�;&�����G=ݯU�����5M�s���q��\�/�L����w���������p��No��6�~c��A1[� �Z����rg��d��8���D�蹣��*����+$.�e�}W-Xm��Y)�yʷ�n�S܌1}��g�ͅ�ep�["N\xk,����W֣�e��Hj4�B%o��]����Z��-��,Soh{�U(��y���fi����9衼u&�"��|��j,�?��jY~�bI�<�ji4�Y��_C�p�y?�F�+�4�*}Zq���&)ʐӹ��E��a��/-E�YYI��zT��^rWt�2����b�[%­^_ hx°wy���{���|���C*| `���2-���l_ ��"�z
�"_�� ��Θ�dV|<s#�ꭇ��":��"��$iW|��5&a��8�7$f^�i���]����0���z�@fP�Kx��;���&=�C;�b�CV�\i�aQ�s�7���
��w�%3���We��:���y|"L�Z:�%h6�Y�s���[⭠��q��>��A�Pmz�A�c�.�[Z�[d��i��e�Lh��pc����h|kZf>",;>0�J���?��Ja,��Mod��W��C��W]�D[Ò�{��&����+y�mUUī,�U�m�o�Q9[�~��沺Ը�n�1p|D�R�U���m� Ü ��t�C]-���q�q�k������r5y�a�87�Y��q�WA֔L��r^%�"�ĶN�w�>5��J��x�t�c<��^���3�"�L���\��R�S�ę�v���6$!y�����>K�(�M�bC�:�|g���V���֣�w��!, �M�mھ��ZO1��w�K���Hբ�˼����׊J�բo���i�қp,�>fl�/�Ѽ9t�?j���?"�޷qn�k���	)�\9�8<��L\�_dr&�B����m�k���l6x����[��ə�<�,_�R2�7��CՇ�vL���/W��h0�J]�����T� M9�R�+�?���C��Oy�K�����¬���\���p`)A+����ͥ�F	����%f!^j6<����j�:dn�k�Tg��5�V�>np[�Z�w͵ɯ��%:�N���z�-�z�me�#��z�f�<�N�Ϯ��yJ�41�py3d�i����'r�q��?���s�9)��a�[�A}7�%�.�'�YZo6e>��[�*!�k�,OwoR�_S��8��0j^8?s]e��K��m�m:b���.�sC��*�FM+h���}N�yp��/�@��-����QFK.����k^?���2\iڿ�i�|F�*�dDE睼�S����t���h�K�?Z>�N^���ă+r��A}Gî�����±�f���P^;Qu��l+ f�w���i���h;�����of�xM{~�W�O��YG j���D�ͷS9x���$y��@E�gXlS�6��)���ӷ�xD^���u�z�D�nK���hҒ�ܸ���^S��g������Acp֠�/\!�pM���G��/��>;�i�:��jj�7;[��!*�����tآz�%z~��Q�jjWq�u&��'ҫ����O����>tM�*ƛP��;5���x��7�����ws���-7�GQ �׿^��筆�����rA$��\c!o�Sςs�պ���a'�c�;f�}V���]��u�|r�ѫ���=�e����7V!)�S~q��I4a�B��Y-T����P�2o<8_�	a嚪�+��4O}�ஂ
m1m�P���b�T�����~4#}��7�gP� T�8�)�� :%,�8�����1�f���8��s�]}hܑϑ����erU�F9�@�s�"g��+��M��n����A�3�6�6-�?ڃ/5�gd��/-1�>��*n �:�W��-�9WҜSM��ț�xg��Z~���>�]>�;[[Z}i)f�s� �BcS�HVӻ��=�W�tQf�"Nͫ=�ǫT����L[�2�|�$�8�Vڧ,�a�,��	˷[��2���J0�&"�ƪ/*wtm�%!����@ITc����=�Ү�z�*�0r�Υ4Bܢ�6k�#��G���i�>r4�]!��5wD"qq��Lk�D��Լ�NrW�J��"��M�7�PA,dD���ZT/����9��%C��s����6�'0�7����I?��k�z"[��a�ʲy��72��p���z+=v�����K�V튫���XU#��+�M�}܍Nj4S*���[EŎ�:9S)t�����"d�n.-���t����/�i\o�h�n���*C�f���r��2���TyB^0�w���y5�`t����U�����+���<��n8�K������R��WI����d�9�B�v�.��r�ލ;*���rh���&�(Wc�%^7/ظ�-K�j��$����b\ދ�gd��7d�V�/���.'҄�_��}��{��s�y�kL���a�"���w[���t4��,h�B�*��`Lb��:w�0��^��Hr���6Q�GxMUr Wk/�7G�e�K1�^����4�jA����;e@���u͘��8*�ݺ4��ǂZ�[g��^��oe4��Zn���>��Z�l�S�X���3y%�ŷ������[}���륏ҖS�&�渤v���3&2�Y�������u4�vq	{�A��I���y�� ��<|n�1��E�<r��d&ދUa�x�'�Q�n�����4� ᣩ|��b�����W�K/����xN���O�e��vBb�rC
�sPB�V�#��~*�⺎#k��^R6������҉���	"�q��ٚ�o�$s�r��q?�M^�Ť9�Fe���hs�è>��
8Dc"�d4��DX����R���X�k?��-q{�|N��r����4��*52Y-�� �^�p�.�^vd.bF���͠�3m��Z��������7�)Z�Z���b5j�v/��X��~z��ҏ��ơF��&Є�W�c���g���瀱ޢqI��z�E��ˀ��\|�ƀ�OrY���ꑯ�O,�����8�}�^��f$P���(�G��)����b�e>(H1�Z����&Y��(`�n���W���l:_`Hj�_5[!��GX�_���̐+�e���?~]��y����Kҵ:�h��}���I|����L�L��pr�w�u�ƣ��M���sWH~S��s���J�9�LB��ϗ.�Y�K�_ �6X�Н��c2���Q�JVr�E���0���P;��X���fS�W�\����0���5��{�z�ד��Z۵j-�|
��7��3��PPq�5(#��h��	JG�8י�'��m�/��O�=m��`Ur��W\�E����C�[=�]��kry�Z��+�{�����Pӽ����l���z1��4��&F����;�[ÐJ|�Z1�D���檳����j�����XLF�(��8�8吀�t��p���sA_GG���Wp�¨�Қ-��tG�<�ZA��L>;��,�R�>����Ą�:��^�Ӌ6��%�!��%�-7���3c�0e��+Ցgx�-�����0��8�.�2h�8��#���AĐ��s��$<l9?��Ok#� �H�ׂ���� H���XK�q
�_	X!K;Gr5���-cbO��PI7+������=���k�>n�g>x�y�sC�13+z�n�-�}o�F����3�{*?�l#𤨡X�'���Z��iD�Ic��,���ž�-[���|���ܓ5�[M���0\��lAme�q��+��!:�ɮ�I�.��<Q������IE�U����A�؇1[�|��&��[��d^o��[X^rs�sBe�wfn����m�e�S.�hEQ>������g�M�z�i�e6���OV�)�|ڣ
��>�#�V$�=�8�CK�1��_��c���^q��@2M��%�=�}j�ġ�tٖG����⡼?�%��i{~���c���IH�~��_���3DO�3jI��E{�.��	����DB�p�x�4gG~�=i�{h��k�l��nÀwn#����$$$�|2��V�*A�oJ�Y�&��[?y��-��)�H��k��˥��'a�����\�wZ~����L�_A�Fq
G��l����^÷�r�/��&p�F��0n���:gBS��v2`�*�T���rl3�9��z>`@�m�iG�}���sFָ���w�ݸ�ܻ���+��wqmw�a|Z���أ��۫$$���W:�G�>7 ���¹G��7;�^�+Uz�H`��C����6�
2����!��Ki)�R���.x�wX����W�P�N?T������31�����S���VO���3��M�.�cw�@y�Q�YR��'v̘�� �� ����
�A���fGO�^���1'>l1�ϖf�X�s�jw��Jb,ELw�����j�g1��oф�[�Y���D+����Eb���-��w���6�����MKߟR������=�#ƥ��@�!��:԰���[n� �����Ņ!���� �C���{} �$���&�r6�[�K��cv�A֮վ��V�����/�����P��s�vRlV����ek�(�v�_b���]����}�#N�q�|���?7.���3� =�U�Y����僘$�}(�Я.��_�#?�Z§5����ķ�⯴�p�!G|������炯�����6�H5��]hW����P�-8n����!1\}�6<l�0�g�5Q�'�x������n�\c�����k*O/�Ӌ������u���m�s�<�ఋ{/͡�C�)�v���Y)�$n����w��<:�P]LU��&�z�:�?�=`�9߳�ab�n��㣑G�u��b׉�b�'� P�w?�a�`��3��]���Rgj�(��W�6�W$ w���}�)�ꊪ5|9��/IMm��g��	x݆0F:�ZSNdmr]��Z�a18@[�����߰�dlP ����T��.i�>���,}��;?70�/-���E�	r���׿?�H�_w�^^� v܄�����D�����P~_9֧�Q��e|"���D ��4�/�2����L�yJ���&�F9����	h)U�<ی"D�e�I͝i��ح ܬ���L~1�I=<�`X���ކ7 ��;%>u��=��3��̭{�����1�J�Eb�(f �葙�/��3L) �I�&��N�N�ŭ�/����X4k4�7�	��ž�2!�'"-�=��O��\����h��P�!�	O�A�w	����Ă�+���a�Fb	q������ �(���-$[n�.8�ʣ.ob|?��K�;�X��������o����p5�?΢�m�l���W��I�T4�A�Su�Ӛ�a6�q��L\�32�� �O��ӈ}�IZ{��I�TB���)���ٰ�*Ъ�{���\�Jxz��?[n6[Èp�"Sƭ�7>]�H���u�X"�� �F
�DGfD���&��2����R ��������I���:����:L���on��*}���X���*-����͢n{jm���x�{�ZY�����ޚ��B8Gu1dҌ���D~)h���8����\�ZL�U$n����W�K���.��lD��*4W�,�>��QM3Z���^�������tFf{�|>�XI�-֞�7De�����罉 @�r/��ؗ�V/h��qs�5eޚ�^۔��!�I�4�̐��~��b5���F�9�y'�2�z�5��;M��a6L��s��h������︎���o.��b�"�]��ĵVӣ�����cH�+���]�&�.�����-�}��ޖ+�U�U{/��N���7�vOE��ɜ��O���]�i9K��9*aٕ��[!��S��!�����<
M����r8s�a/SCK�K�u D�fq�	l���Fe]w.s"�
�-3�\��0�$�M��|,V��a��	��t��0(B6FKi��Pҩv~FU=�r�3��kZ�)?��|�FM�@�۟���nM��h����.�ۮ[��.���%0�u�#XWa9�����wk�
h4Jj��UI���Wj����uZTҦ��\�z�עO��N.��)�h �!�Kp[��aV�]E����z���^rfl�^��[��3������R=@��{^݂&
aސ�!0Le�^�c�����1��I��pHq쯄�����]wD�2�#���ٶf3��������0Q�b��Rz��+����!����{��o�"8G&Uou�j\�5��}�$^v��W�|:$���j)0}�[VW�����#\�}�{c���e"��ẑ���}I>W3��c��Հ]�0ߍE_"��޾3���>������c��v�!�7��T�wV|�"x��t�B�ٍ�0i����#����åXIr-%��x��{Ev]��i��C�>�-Q>����\� ���i�݉�կ��!F�r�����⤑���;�{޸c�Y����#&�Q�*��0��y���4�b%�p ����D�:O}^��VE[1�P��I�c���B-D�>Qp	��μ�[�H�VA�D�7�bN�b��=[�����F��:^�^l�#G����3\�WwU��+���7.��Ԉx�/��>y&�m�E�I����/�n����&�$G�����'vB�3�<R�b��s�/� �G��&��;�ka_�]�N��܅�ҳ�B�)C3
H$7�QCV�����@���*c��� jq�7Wx��T��6 } �K�~':�D�[���X0���[:��4#�5R��ɻ������٣�V�9*�R�gؽ��?�6F63?=$��	67�b �C�"�e�Ѻ�ܹ͐�?9�Lf����� D��R_k��.�S�;K?H5DSiZ���us����U|8񁖨�B��M��c��&�Tnf���Ƿ�D�	�������U0�-?��?��6�g:����&��6�\w�������봉����%�7|`�'��J�≩#ĶNNHK�xɅ��_h�Lմz��Ņo��SW8>$����2C�ijjV�qN �$(L4�7o�eK�X�' CW�^lQ�7�H!��)�@�Xg��{����d�YR{}���f){��*���LtA:�#R�V2
��>��jY����`�B�q�������3}y���9y�����X�UcF&�c�NY�JvF����?�,��v��6F)��g�q5� xP�&��cƘ��gO��W�2&!Fs�!w[w Z���K}���5t�*D��M��Uc>���� �z�S,cb4�:)�ܱ[w��^W����,D���T�F�}�x����b��"�¿�FSV���b )+XAu���0�34j?�x/�&�Ր#��H ��^��ATұs�J�0�E�+�j�ں�;ֱ����ᅅkEe�咣c�&�ƫU8�r���y�+ NJ���Fd�����qx�:���g+��e��s����l�ǡZ�[v���?��dbYXRY��?�K�R=���<���pV���OSk=k����`��4�����h�5�LBB��͌
�}��������=<���-�:`����H������!��g��_{���s�(���̏�����?}�G��轢�y�UJ�����l��D���Ò[��W��7�ޥT�omTJ����%K}b`Μ(��^w&!O'h��#C�޳��(���F���I0��eqex5-���E���K���1!�F$�Y�Pi�_�R}� {�/g4�l���j�zX�_˻�N%��8����8��Q��g[�5�W����jJ��V
��A�z#gEP�	��ܼ�oLh�,YQ�+d��r%nv}�d,��@Hrz*:��2�' ���}�b7P��|�NLh]=�s���'j�X|��녾�B��NZ� X�[��W���8�SQ<�a][��8w�J	8媿|��6\Ч���ͺ0�B�,�e�����]�=Oh����&%^2�Ɇ���@�w��DXmčWU��}�oS��j�E��S�u�W���d߈
]��<����c��ݣoץ���ʢ��\�=��1z��I�uSŰ�r�m���/>��O�m��hW_E[%'Lt-��լ�z�Ԫ2����/�^pΤs߼qf�z��r�|N�R����ƫ�d_��L��jkg߇,��Z���Dߨ����ڢ����O�� ��i-o�Uo�a���g�~ϩf���P2f�����PSY�#��d��:�,w���G�.`� yY�{j�6mz�a�K��s�AM��йZ
# �~I�-4hD����q𘛏[�4��V��,���x�߮)�(��
����uC���D�GA
����`����T&�M�"�bvP65�=�q�Z^�lh�dE��*Jy~>yB4��;�҆����;��0~Փs��h,��7 v��|�uK�՘����^�x�����A�����=w��)�[zs��Gǥ�GZ�2FЧ�?�i�й�L��9�  M|�P�G���<���{o5!��&j=ڽ�~u����>��F�5[׋ن6ޘ��ʛ��A��d���,�@�8������Z���z�/�U���9k���y�j^�<B��z� �s@�u�gf��}�K_�jE��<���7��˲ju�wC���4�b�����B��&=�A?��;��-�)��S�7<��/a=�R�iIAv���.p�nZe֓H�GNh����AB�w������a�|�/HI?��︀�� �Q{��|�ۢ�i��jE6x��4�ܼ�]�^��8����Q����Za�g�q��j���PMf��节�(��m��oKKF.2B����^�0~��Y�$,�}��s��:�3׽���X\��sG�eG�w�ؖ�w ,د����گ�]BȈ�"o�P%oR�/���{��| ���$� �����m�f�a�dՖ�O]~_%�	�n�t����?Cu��?�9B�93я���d�Le�S�te6�sֱ�ܼ���R��=���"8��̌�@�q�'�1�5@���@^:�GX��rt]oil�9���L]S��-��)z���{�L�ԯ��%3���<+5�"yӟR�5��������N�XַJ�}���YM$�.�kE���z�1 #.��;�����*�A�Z�ΆY���S��e�Lw�;����4�9�:�Ư^���7�ǀ�|^X��#�D�	\AKC�h�Y����1��L�|Z�����l�Yc����ԃĥ$��]�P2x��H�,���?Zu�_XGT�^/M�?���u3�4�3�v��:X�EM �lm���P��^>�o%Ϣ����5��	�y�� �&��+�}|xd$�<�W|��������=��v�:ƹ��a���R󬝃:"ѡ����q`E��:ƹً��iX~1rgj�{�c�2���� �쯭���%�ò�>,a�&�A�k��8#��u�z�x��4�k*j�7{���z�9���>�	�#�`�G��Y|�=�j}��d�BS�$j/�S�0�q��'��y�8\�nLIEs�<�۩��f���;y�H��#��:lQg&�+�l�sϭ���bÛn��W �t:Ƒa���2G�Zh Ũѹ��KV���N�6��$`�z����ƒ��˖ ����.XE7�L�AI��%�	�>�+���~�-�[V�~����������kP�f$�����Pi�����gqZ�F��ٽ(�lH�8�L�}��ٲ�3�/�H��(�Qzn���9:?@3%�W�<�����<7��I5}s+���	�l�����;��;��aɢ@�T��ߎcU��uUkuc"��K*u��+�i��aA��)N�V���~��E��2�\i�>��́��s�pׅ�渎y����AN��}���@��*�D�6�A&�!j��*
��T�;Y,=	�o�zTY[���N��گ`��+zt�=�6�ia1�?u1�I¹�����k�!�$�d��2�ɠp�tZ�8U���ySd_ ��}H˄�%��<��H'���qk
�-n� =�
k�'h�t�T+��v"Y(WKZ���P~p�S�JE�75��ʧ�Q{�p�� �B�Lm�Fw�.�f7���	2C��;���	�x�	�����jJ-|vcz��<7*'��i�-�ʪV3�J?fFJ�b3�/A�^�B.\��EV�xv�5իV��{�9]�C�5=�-��ּE,����q�ƥ������M�Z��tY:zu��G�XĻ3o�	�/��
|y ����$��-"��ɊXӝZ�׼h�U��aN���:)h�e�ܭ��fo��>:rp��تj�([.jsD󂗽�9T�/��`��V�6����MƉ٥�MQP����q)]wVD=���)�5vFI�e�	0�l�}��^]`B�ds���I0����g7.�I�c7u�bTҫ&�GO������f�P���lp��ՈS+z��p�ys�a�b�`6��M߮�L����/*� ^I��l�[���a�"(�)�v�\,�z��!�A���5�$�G����"�7~��X� q�J��\����ݟ�٠קfyr.�����KM�S���e!S�g}�O�2jJj��d��{,����rDK�'Yx��IO�QS{�u��A'��C����z*��$��N�u�q�+>��@hX ���[|S*Fz�iŋu�l,Q��q,^;ɰ�I��W�R�����J\��U_�/�A���!��PRx�nhF^���m��dd7���60���M�����UK��r�:��t����rDK�J��Y<_����J� Jp����W
�|��6d��
�(P�Z��]��=��ԎN�BN���Zм�h�8�h��w� P�����v
����e���q�J�-]D�������)�,���!�9[!?�yh�=�l��U�UK���<g�@&p"&!n���z��L�j%�u,��5G�7	|�'1��10: J�n�0�0�6j,��O������&��|0h�sG����s>N��
����kW`�6���b����iHL&���.tK-�i�ƃ��(3� �t�۽�����t��m]�ɀ��i�$U,2��h�U��@�\A������-׶��}�[�d� �x�2�v�>4�ysr[L����S�v�⇈���b
G�I݄�p�r����BhnJ�H�5���ic������,��,U��{�O��[��N��Y��.��Á�@���5� �����Y}��K��p����w_B�"���5&��v�k��v��& �O�ڪ�k��س���Bw?14���.��=�.��&x	��kFf��o6q��"�=b[�O��ۿ4m�9;���p�}�j�[X����Q:W�r���~_�nw��F:�l_#�����<�m~yy4�O X �ϔ��|>wg��iy���C'�[�RM�/�F�QF@��W�ܵe�^_�ih�:�ݼ4��q��Z�C-���Ĩ��`�TYDN�����ʡ�GkvϜ.db��&�._�P<��ۿ����N}�[Z�%��_�k&�u���v�\�_=Ǔ�S������ֵ�J:�pz���/4���z!�
\����{������e��J�R���v�KVuw*�>�Ռ��>y�_Qm�c�>Gr�b�a�T��x��T&���.i�&����� ��c��^�oe�ozDrg�H���0����H��Q��	�z��� ���T&�u��we��o��xHn�WF�'�����@���R�׀��b�oʗKg����6��V�wBd����;$��	{�����ɫ��b�~�:WȺ'Ə�g�>��Izއ^�cK����%:NǦe���R]Q��C���uǴE`��6��H)*�Cw]����?��5�~�]�屧Y�T���;�8p���ull�%�S�W:g$���L��:�٣|2����>����
��/��p&��������\�_T>�4z���Fҥ�w�O�x����ˏ*K�f�%�\ŏj�OV�k�e���U݅�f��y��)cЦZ�\�nu���ߎˁDʶ����?43Ph9 �+�����@Y^�gP������샭}�k�L��ħ4~�qԠM�����[�d���W��AH�R�~�o�y����j6`~cr�)���1y��<����Аx��)^��=�`����[+��Y}���-;x@�g���*����T0/��[x��9 g��{��4�>�K2�\�D\�[�����K��P�Z�j��A��~�ć��1;R#��S�wⴞ:߲��5u���M�sʶ�������r8����s�B��*��Y���.� Z����C�ȍI�@���uV�/���Y�=��8�ˈV	���p�, ǹ���i��G�B��W�������j؋��
�WR�j֓C(��x�U�)��0˻Ƀ��M�������Ӄ�lo�g%�sG?��٤���j���'秆��h۷���ŭW2aUT��c�Ñ��}�r����ǭ� ,�?��q�C!H��D��*��,�u��P�p����Fv�@�}�����C�����XV�]�[?�|j����rA�og)4k�^�ϑ_�Wr�y�]	�n���;g�ď{��?���o�#�����Ϭױ*'�;~��ֹ}�X>~1ޅ��
(��y&?�A$�ī�����wȃ��z�Jn���9#�e���B?^�6yS§޷"~n��b?�h{�e �&��>�3s oDc�BR�*�,t�R��fs�������3hF�	� �%�l�4�@��z�{iԓ��"��3�lpF��8����}]���- v>�(��a��c���D}���W\�ҙ�N� ,�H��>�i��)�S���Զ(��9��:���/v�!�a4��$D����U�7���ёCdx��O2�
��b�ĥD����1~h�]�����lFd�#��i~����r-C��7�`�c1o�ٹGNi��<C�bQ+��.������9�D�(��3���Z��H酘��	��e���q�aj����Lv��u4�6�:a��/��g޽�>)������&�/{���K{��wu��Y[�Z���5�Ƭ�.+�G�ݽy����"����ձ�b���y*/�T�)����U�ϟ+8��-���`����{ƒw�o�sl���s� �d�����\.���ÿ�A���}=��[�!=�L��R(i}�����L�C^�:J��e�g�D���0�߻�H�i,�S(�Og�sV��"��j���P�~yj��.@�"s�Q���|�R���zi�&`@��*����]
�7(�k.~~���m�t�v���ї+���9�����,�%1�)���h����A�]WL�Y�s��|o�)_�i��3����M��Ƽ[5>(K9� ��X��������A6���>�%��	}mUF��Ah��\��Æ|Z��0���Nwb�w��1�`��i)[y����7
����4N*n�Gӣ���^�-Okdv{���|Y����2��z�r�؏J������p��ZP��������W�?��M?p&`@dc&-(��G
±C2
�P��$���ju��3�M$S2��|�ߪ�񿒳"�a�D��1��>���_	�m-Ş��!�_Z�<;��a��t�����땟/iTQ��p�Pl�ݝ*�E����qޢm�&BR�#�����(���E׶�G��rl1JQݭc	�ڞ  w4�Tr���1;��0$s^���CKv#^�ᰕl��7q���F:�����?�9z�Eή�����t:���[��*U�H�M�}��5� �gj\T/��߾l�����[�Y��:���t����&|����-Q�����a��uHh����9)89�����~�5�_���휝���Q�xI�����6����r��h���2B����״�;�T��;�(�DMޮh%�50g7P\CBE���~ݪ%�-��Ⱦ%����� <���U��7�_���_���yU���\��C�?�O���m��tq.��_��v_I���fw\�U��MȜM�޴)h2�|�&��"X�V%��_����3�"=zN%z%��U���⵼g�Fۂ_��g�=�v�8��Ox���F(���W��qt����.7r��H#L�YF�*�>V�/�vpR����<����Q4"�;]�"�=�|	,qA��O�i�9��4�É�q�V&��$$ɷ�R�@�j�c����(��x�]����m�U��ݓ����]ܝ�-ʥ؎��>la��V���7/L�ſ<���x:kM���������)j �@�ԣ�AU�?[��T��ne�՚δ��`���F66��O���s@ם�PZ��E�M��l��:Gd����!\�_����6�	n����j
��n��A~
N�}�Q��KuPOEP��6��ę-���V������>�^J����4z����Wǅ��\KG�qq�6T��5�ZR4υ<�o��o}��iЕ�0=ԃ�b����O�ǏkJ+��n���G����)�c|������.��Ӵ_-�*���!�M��G�n�*gO[Ɠ|$�6�5W���qX���R�!{�sS�6��ÿ��OWf/��?S|Q��a�G�A%���a0<A�N�g��k������}���5ۿgcWy}�-_�P�Z��`7�?u6�m�P��B�.��ƞ5x���	kn��/�M��,"���9���?�J���%O�(���n�U�B��cWcͿ������i��Lm8�\C0\�<u��O"Ì��P�����0�+�������j:tZȚ ��}t�ьң|9���k5���-^#�����[��P�K����x�o#���^vV�/�ӮK'�0���+���2&�TSKl�T��ԍ�|ґ�]գ���^�����N �p�	�ŋT������p��]%�a�v���q�u��%t��Ƴz4k~]��L�d�ҿ][agscSԩ���L��}�B���X������R���)�^��=6z�=���.�v����IZ��B(X���䎷�ԅo��4�<?O�|����ٛ^Z�/>�ܲ�_^�3(}�Z]x�Y�k�0�^�J���2��&hz6�p̈́&�����|��qw���͏���_�Z�H���M��[U�|��d�kk�ڊ���LU�E����5j|+Q�}�|+<���G�]��	�MĮ7r�FK�� ���o�OF�6�j���w�,���^�1���x�t~{�W^1h-�I�[P�H��_0þ��*p��뢀KL��s���zQ-������;�Ml�&R:��Ǫ s�
bf,Gf�uv��#�����^=�Y��,�'a_ȉ>Զ�Hy���X5��r�޽�W}��l��9�n������6M���q�0��~z����mny�ٯ����q�4�0�7���ު	!/��.��6DۓZ@<�UF�=?�H�VI<�X����^8�"��}
K�j�A���M_mo�ZL#-����j���31��o�Z�A���"�v��;�}���y~5b�~��_�1�rR�CN0��˛]͢���̠�/s���P�y�X�v�%���z(��=ԪsO|�y!PV� ]�ES;���ޕ�F�z��TEj��%C���ߦ~�i�T�G�-��c&�ҵ�w(
UL�?	i�d��Τ>��y_+h����+����������[�G�+�0����Z�U������F5�$�����l<� }q�Lm�����fTR�pӑ�3lo�ҩD�����=`d�١X�;�q��(� ���`TXÍu�-�LS~#�m�����Yu�Z��>І����^���QT��=�d������}�R"��GԞo���6����������2OvS)\~��^|�Yp /e�� @]ƹ3��� �o��~,Q��l�`ӝ�ː�Մ<��ǿ�@u*W�n����L�q�����J��U��c�Xq�WѴ���0�ޒ�{�l��Id��oZ%5y��ߎ�K&$v�V~	V��j��=6�@��n�y���ۯr�|���~�*Y_�L�^�(/Z@j[��TT\��3[���̮���Δ��Z��ڮ��L��<�@���˚�h�jUޙ;��f��$D6���f�ié4��"+$�>��B7r�rD�p54�vB��_�u!t�h��&#��S/�2BH=M�6�7����db@-Z]��.O8Ҷ_j���,�v�ᷭ�ҞG$��x��Z��`�w�.���q �����˹�f0X�?��z��ͭ�Ǿ[7��}a�5J��.��݋�Vp(��^(n)P�݊��[���	�����g�?�3��3�!D��{��>��I��c)q1ee���������g�E{W�h]k��3�FRs�c6��MNj�\��|?������ek��,�)ru�[��P=�Q�
*�9@P����8޶�����WɊl���\��/w�b�1"<>������#.����b>��r�,hš� 
�t��W�&D~>;.�C��A�J{@���?�7*S����~v]�m)��t+�Vg���-5Q8��Fw���7�;j]q�"-�#b�����"�5B��p1���;�/sF��`� f<ܲ����8�H�	sma(�좳;����>\�x�9�5(�da-"��⎡��_U�D*��^�0 ����L�E(4�=/{N� �����$9��t�
"��8P�o�K��pW��N$00U� ��s%��|�Z�)�م��,�KF�T���I%����ݥl�X2��D�^m~ˤ�K�v����@��I;�Ґ���@j3��FUj�(L�Y:�)�N��
(y�qۑx��G�s d���O� ���(�HG���B�s�7�L�R�� ̉�2�9xE\�l�`;p>���
(�I�7�d9��ۅ��N�&s��T Nx�*q""̙}���뚶�8)�xg�I��r��k&���(�֌�1�qd�.��DEK��+��^_z	�y��)��@��um�|�U�R��!.����Y#no~R09�i��N�Z6mJ;��`�F{�RВ"O����Mmp�Ia�,��޴1�C#�|z�1�ʭ�Gy�2�H,�����tr(D�WK������!]�r�X4����V!��(|��SHR��E�����Ǥ�B�:��(K�Z��S�Z�<W�c�~�j�]ڍ͠��[nΈ�>�UBv���-ݨ�N����_�6�R��Y���⻌�R��e�6�@���s�B��#�Z��*7�����|0V8;<�ϙ���[��EN�6���ߝmd`�=�����W��e��O ӱ��V#�ĉ	��}�)�	�{�7�e�``n�x(=Is�#��Z��i�(M&g�����oO��e?��C��V2��RyW����<j�nL�C,���W�G��=�3 Fۮ���v�/�޸ �a�I�0
6�`1w4�q��R�\IT*��y׶�*���"��H�Mᡛ��̷��byAϚ��!�[i:�p��;D��w(Ć��M�/isK�[�ˠ:�xS���)iI�m�5�c��©�W$�A��S�҂��Rh3�Z���}0,7y�w\,J�R�3���'�PB	���:��7��@<&�A�!��D `G�d�(|5���׷��Xr���F���RId�iڹ�v@����*q��X�����[r|�����+T%�X ���&�E�f�+��a���G��R�c�D ��?����qp**���� "_�4���n����i�����ǡ?1ˈy���|)8����$���(2��~��da���m,%��Z���Lk�m�Q6��)�-��lWM̄��C;k���x�.w9��ᬕ[ߍ�>������C��PY,ݪ|� Mi��y�x(s���e&\����9J*Os�����/�}����r, tadmu|:���y��RU=2��SM�q�_���۾�k>9
ع*:���@�����g���I�'��U���%�+H�~��/rr�G�I�u�%W/�������J�Y��"K��4�(
s5��ù=�t}5�N����4zW�����ݣp`��Q�Wl��H7��ys�����&�^����7=ܕ�d�.�Q�$�G�Μ9� @�~ q���[��h2g���h��=#��H>��Ѵ��Jq(d���H�:G�WV�3�Pq��+���٫�� �S��,z�`�V���(��9U�ߌ:�����W<		NX��E�����)J��B(�YJ�ݘ�F�V��q�K�2��! �N2.1J�Y�QB��$/�s���}��M�\ߗDi5�6 ^�S�ɡ0 �H�_S�p����C��Çi���-H��|@1��!��j�7�d,>�t�L7��Dq��lp"UuN��S�4c-�bBWs���>�JS���a+.dcJ�N�9|�hn̛���ɧ���_B�7�+F���Oz,0�b� ����r�Wy�Y3��t��5Sia�me����NqEb*V5T'}���"�7���M]9b� ����~��-[��T`x�����W�{�_��_ȑ�\!v�*S��Oa��p���3���C��M�j(���Y���٦U̗s^Xt;.2u�/�����L	S m��6����
�m�u��4�z�b\��{	gDz������O:�M�҉LH���C
$�|%g��Jn1���O *���J�o�cHo��ҏ}p^����J��6qh�7}��]�[��fZ3t��º�j��r�� Z"ӻ��%��!_�8�8�d���V��h �zF�هj��sڗ	;|`{4����kh8�P(�袙��ix�K�x��!��[�������OW�»�5EX�����XW���X��C�0�֖�уSN�W�S>@WR���M���F�X����.��7�XN�и�>�v؅��\x��4S��ݏZ���R������)���\��6E�:���j��ti��q��G�'�r(X�y�\����)0�D�Y�1| �Ȁ\��s��}�<��|��8b��3,Ɵ�k<��u�2^k��|6#�րL�Nr����I�tj�T�e�k�A��h�#=U���7L=���VI���|LPNo+��	���o!ۄ;HU�h�z�)�*d���Yd�X�D���YJe��rN��I��X��]@�y���	
�n%!��!�kU����Y�E��L��4Q�󉾤!u,�{�4F�i��ly��"�n����pOv�ci �p��3#;�����+������e�3�Q����)�}��o�r:妼���������Q�lھ:zWr3#�p���f.�_%�	N�\5��ߪ����MgW��F�\�c.� ��O ε��gZ��u���W#~4/7�q�m��u��^�+�d?Ne��0	�X=ҺrǓ�?E�q(�S@��������=<L; �:��ݫ5�����Zy����Ŗ9`ɛu<|�~M+��.eǾ���g�k�է��o�S�{u�j�g�
B���)[��5��
�,[�[*a��L
���F[I�h�G�~߰4(D�N�RȨ��s^ɒ�!��V��Wz
�՚�dI���2xE�~�[���YjL4i�H.:D�S����s��t�:�3�h�����"�	�\�$���Zu�����P��IaXhAt\2_OZ��d�:U��a�tF�DkƗ�'��졫�݀�������qi�v�q�ǵhLbp	>���a	���{� �ty ��}z��%�a��-0��AO�z���L�Y+�����H�7������ƨ�\4����1�����p_Y\?HH`Q^rH���H�H�����pO�>�o�VY�i�� ��������0$���m	p"T��X��'F�Z�� �1h\[��|������P�B�~�0�$�n'�px|�X?re.lE u�ё�̈�?%.���� ����wrׇB���ly]+T��V�v^etmI�P���1z�Y2 �Xc<o ����ܦ�:R�.f5D�`�b^�g�xL��Eno�K�[�"����mRH�OLT�_Gi̊T6�{+�h\?���-}u	K�9�a@Q2�1k� �J �!���K �ql=s01)���:��L+uOQ>_e����?8mNpB��H���w<A�����{����RXIsA[�V��w\ȠC�r�rC��;�[���a�h��؋*~�k��"Km���%�_v"b��'�0��#Vce:]6~���0�`���]Y������H�3�Y���idk�j9��e3�)���<��ӹ)�^S���������/U��2��vZZ��k���v�t�M Y�ȉ.�� �Cf���Mg+3r��w��9@i�֚�q���Ń�HaU������Qde�>ֵ ���z�*�a��F��?�m�q�)�̲�J�%�a7���9!��A��9��x �g���!d��^��jN��faKtn�߇p�y	�O�$���!�e��R|��[�-+AJ;WE�yƴ�=G�K)��/U�I��5���pZ:��]:��T�* �� �V����3�߁�s*yb��J˜4�7Ъ�yX�?9ުD���e���g7������;w��p r9��ʿ�y�i��f'��2#��d�
=C.��V����j��(�
xt7����r��&܆x��_������X�� ���Kٵ�r�c�R�|Z͙��CF]�FO��~ ��S/������z�SM�e%��@���]�:Ŷ��gY�{�o@"z�� ��3�+D�K����%�8�u+Z��\�(%�Б�ðr'��kjd���.^���@�\`�!!�y͓I4{���)��پ5(βs5X�k�=��Ֆ����G7���@���r��c�9fa>�Ek�!��/V�z�&Sk�C��6��M��ޙ�W-�~D����s:�=ޗsض@&7:)�f�0֯v�¨>J�c�^���b�+� ��<">v��+��V��p��7sIB���8�� ���T��3f/���0�n#s�BTK�P�$��7���!<�J=c_�Cd"��Yx��6���U
��Z��B�s��:=�t_�?
(q�^�D�>˔_n�tv��� y�	w*�P�<.uM���5%��H�f�?�
H5�F�d���b*�)�R= ���e��� #��{c8���{<���ZP�����^���a<}E�]���!KmGLϼm�XS G
uƣ���7�8�2�,P��N*�
:J�e�Ԁ���
"p˟7P	0�{�/�咎�2zh`倕���{�%����MPت��n��eX���H1IW
P�Ğg��}��)��S�tnp�۾
�|����n� s�b�)�YT � ^
y˥����ߝOR��S��5c�O���d�j�e�/�b*���.r��Y\��J�ǣ\U�)���
�������d4�����4��<�*�Z�/��t	��Њ ZTfq������Wa !�ع��&�+���V_��uo��~���e�Z�8Y"�G[�]����0젢>�Z�+��9��
�����=têW�G���hb[��J� |�6.�cn{Bd2Bժo��}���OL-b8� ���k�|;Wg\f8��/�?�V�����rN���<lpX�)�5T�OQd�ON����9C{a2�J�߷�ut��~%� ���C	$P��(a;��y�D ���I�����]� ��<�����L���Z�oJ�oJ��S���G'%T��ð�4����*�wN�-K��:�z<����Ev����U��e�/���V�HI�-���i��� �r��F�1�+�b#��󔤣MK�����zk;�Q���U#�����l�f/��|LRu���ٿ$�f��q��i�d>jӁ+.L��n�U��f{c>�Wx��j�L��2f��ߢ#����D���;��٦�շ�P�l�ŋ���B��E�+.3����0��Y���wmE���	FW�'���;,m��Xz�o_�WE�<�	/|��i�Y�M�Ɓ���͟I�w��<ܤ�� 7ڃ��-8�@����X��.��|Ÿwn��Ջ#+�5�[����g'������T���Ȋw��Ƹ�m	���E�{]��_�[rۅ�l�_;9M�X��J�u��,U�M���f�o���~����Be�cɞ�f�8�M^�=�҇�
Trr�$�T�/���L|m?���f��^��Z�❮�O��@����h �L�2���*��*Jj��\�2hd�k"��3!-P��g^�m��Z��䟕����)�����%�
:�h/*MOU��l����qs���(WS
Y1� �����f�R�.���-,����U^�����4�$�����i�ɽ�F~B�����*��w�ݱ@� �q��aQVwE�.�r\�D��1��r���v4<������0�r��q���i����=E.�/0<Y�	��W�l�p��n0 ��� ��S�i(?=�?�"��be�|N�_!�q~�c?V}�%���m~�́���?�}"�C ��QS���#�����B�u�!e��߯���|��j_��d��؎�(��6<� @�y��R䩃�W�RD*�x��Ȱj�E���G4B�_��[�ѣ��D�$��E�͚ո�V��������ND���^֨�����H����Z]B��n�Bsd��4=nv����M�U,h�|�/_Nc��U��J���cå|��r��%���m�!��	���׫�����?7�z����v8�������(C�������´��D��]�~h�T�Ƕ�P[n�%�p�p ���2��,X�l��Q��J�*ٵ�c�EUw���,=q��<<�����i􂙏� �U(�0�j��y��Z���Z�n=)Z�쫡���욳�ml���i�.]*s�:|���9�{zᧄ%Z����j���<N��H��*�������V�Ss�(��1��?w6�3~�r��]���F���\v���m�-}��X�a,�+�Z�g����c��&-�6�IR��X�G6���o�ON�0�C�wg%g���,��tp���ő-�k���(��u�HYN����^�򫍤s:�꧷L�▂���MVr^�j'�$���c�a�<�퉥��J�O�D+Z�=g~�t8�n8��͇������@qU[1S�ECu�;�O�㣍�sa`�%;�ʌ�d�;��Ė�)>9R�t���ɑ)J+�\�_ 1AY��y*灱�~��pV�g��33¾�߱��h��Y���C���i7Y���|c̽��-Y�S�A�/��N�^��l{A�6��.L�X�z:[1鞼]�@	6���2� �~g��bP�^P)}�=tm5����o�u9�ȏ������a�Ζ&���"���-�]����1�u�R����Ov��4o�K�@+�/�e^��c����5�2;诅6ӑ�L0kk-+��c�5+N�lSy�����z�z��3�в8%yμZ����o��<?�{|�?EA,@�Ƶ�.Ə8��q0gW݄|�!S�p�B�(�k6A'�0:�4�x_�Ce`�><�d�����ym	X���5��d��H~��٭�>M=���n�����a�8�(��˶����4Z������CT��<9]2�~>�T��w`K����3���u
���!t'�i����7U�'W��7t����f�@�w�1��:u���yEܴ���^|���:Y�a��=�� J��\uX�1�㲶�q$�m.��$��k�`�/���e#�^w}���}`���	�f�W�pG����}������z������?	t��U'�a'"Ȼ8@��Ƅs�7�N��ɞ��������!P]�8=\+��SM��d��)� (v��!�A_KyZm��!�������N{�~���䡥Qg���E`��|�^{�x���� �ͽ�AP��������F+�&��1����[*Rjۜ��=�c�Ιi��C���CCiw�}�e��S���S�)5��.������[�N�v݈���)_��i !�;9B�ciHWf8�4���Ѡh�o~FK��N�.�B��~G�ϧ�[���KGk
�gX��,����8�YAI���BM�44�@򻣝�&b�].Z�#A�`(��H�]���b����t����	��Y���u�s���7y�,F�)�~�%P���[V��E�	r�rp�u�`\�]�<���\H��y��!}:}$����}�@�f.�^�cc���,#�p�'��[�@�֑���c����;M�~&r��?��h�?�q/&�I������ߝ�0��t��i7� *>��'R��wsO�E�d��qz!�����i���vQjv�#@ ��&��:�{�.�2w��~�_]���#GC�������ٷ�vD��g%
I��!���*j�=�ͧ�b�ڒ}1�e.R��J��pi�zX@�	�kZ_���Iwt貛Q�4�R�ܷ�Ыn=ݗ`c�~8)���k��?%.!NoUْ��1���؉|jMB�����������H�y1�\�t�F���D��z:h/����7�ޝwp����K�oƊ�ռ�O����oSΐ�p|�!j��mh�Lj�Đ�h���O:��N􇝻�#��M.�{#@_��q m��ݹ22,}��T�f�8q�H_������~�̀���ylՆ

���0�N�?��5N.	���ƓN �S��-���cx����@�Z˷*X}�S�lL4�F���'�{���-��.��L	��F����Ĥu�:���`�]�	��1����@S%g7�j,�v�t ��V1�����u�����N��������}��������E�ط���'/�>��e@�uc��t���[�g�C��#�}��D%Z�S����6����_����M�|klDvL�"&����r�l�X��G�A~(+{��
��̸|��JZ?�u��o����
�0N��2��RYse�*�@]��O�3TE��2Sj���,Z�~K&����h��6�!&���l8l�G�7��n@	�O@����
�
�0�(p
��P
�N��}��0w��F���5x:�����F�q�x.�:R�E�w0= ���n����y��t��i�����w&�x���0�e���-`�#���%�F�FU�8;��9X[#i{������J��� �:��=�Us�_�7�w���u&V��s�G��@n(�����ak�γ���n��:ko��H΂��:��A��V���F�=��9(IWb����^�-����9����'�_r%O�Eo�X%X��� ���Q�[x���G�� ��|E�λ�SہO�Pt���
���6�����귇��Mȷ��Nklּ{]��-�[�7��#���F*�둼���󱙂��	�����T,��s��.��XG�)�wx���cԑ��n�u�k>�Bւ:�HC��e��X*x�1**�O���u?n>C���W�V�Z��Y����$���M�̫T��^�ހ0�5*��0纁䛁38zQ��G��̨2s�1� �0��_�����V�~w�/��&Q���XSzv��3�eKN.G���H�1l�̺�\�zJ�K��Y��
8Fl|s�g���0��c59�Hm]]��ԛ�c�=��́����@۾�T?E�&�L��mdW{ࣸ���V��8.RpZHf���x�qg.O�Ծ��U�V;Vi5Z A-�� ���@�5��h�j��"	�a��ӕTW�����@�V�i�]�E����>��v��|�/�EZ�~6��퀫�a�~�b�c��~���|E�� �| ������('�`��?�+�:|�&/eWDN����5���d+zx�ui5��^����� �;t���Ud��Ek�=k;Gy��E�mz�������A���q��Km��OW���N@sG)Ka���ũ~��q�㊿��X��$�2g0In%�Ct}�p-EeY8�mt��Ľ8� ���K���&�x>��"#�3���Qw�DW��T��G��ٕ��{M�3��ýFũP���i�	6f�{�~]
ԕ���n^߱
���Yy³�v#���ç��wj�D�xZ�B�X�Ti�kHG�#>���3�xJr������q�0��e��&�����Х'G_a/�]��� �6[�ȝ(�B�\��*�;�Y!����?8��K�<��A�b��J��q�abSE^Zb���u��>��7�����H&乛�T}��z6ݔ���W������#_@NϩǇb}����>Pcz!�^r���N���L���xy�X�lP�@ �f��A�6)LVN&�!ٛ�/gwm�V���3�Jw���3Hm�{�R��Wzvx">��9S��S�2'��r' AXt��?�<�*5;�+X��5>F��*@�����v����&�^ʛ3�j�e��${.�F�:f���.g*<��V��N����A��2ڬ�s����K���'�"����Y��!e��+k`Α�����Н�E�V�ܶC�e�(M��|�0�%��?���P�y��dS��s{�G]I��b�@?wH�)����:��-����g�#��Ӵ/6�����NB�u�oۥ^�L �������7��K/����EP��뻇��O+S�q�
�4��\7���c�U�k��fIx���yM�M�����i����9��������v!ֹ��S����^��:���"ZP�Z��j��廞������ڽx�&��uq�� �����������cb�t�!^'����T�itC���59�L�-���v����Gr���Jf�n�nV�2��>߼}�/%]����,��Gdj�f��m��X!xX��\��� B
���\r*���j�� Y*���ȉ�����[���j��u�5��_��~0ً��_�
L+AP�=d� 5#㽳vk�V;c��5��h'wK���^����]���m�nk� g������q��NT/�ܱ[��E����e9���<'��e$)UgL���Fa{�����v�H)o
��h���yNK5n�h���[L�~���ʱ=} ��F,�����Y�he��[�)JW��|���Z�}r�y؋dH0"�}����Q�!�vA�o"��Yt� ����d�~bk��Q� �E  7��c�{����;�"G8�^�9�q}��Pmz�G����[��B��$�$X�k���h���|��V�~m,��T^-5�i3�߽�[���?�P�#R��^�(zu/�>e�Ŷ.��`���"f����8p�ǺO�d��>ϱ�8���/���ov�|>c4F�0)��s��e�v�4г�ɟ|�t����h����7,�����p�����3����U^�n��=�ݯ���Z��νm�ޗ�>��?Eӭ�gtx��B;*I@v�Q�A�+?2*���)�+��P����V[wS�M�*�<��B
��r�}eM�͒V\�9�/�#I��˔'�6ۯ�#�7x�؟�L���$w�D"g<����ԁ�ɛ���a������gM���y�&�}8���o�.9� rZ��ӼW,�?�Ē*�����i��� A_���V��ݭ#r�A.��4V��s���B��HC��僡E �i�g������`m?W&��������Rdu�#����}����=DY%��N��|cA��^�7�N-����KGHJtƧ����{�	�/��L{h4����)h�g,�̀ja�w�%&����5;`��Bs�u���lE����zehF��?����������)��:.t�/D�w_��5?O�#44p�vC�\��{*�8���u�D����k��c�Q|���]�-qfS���""��1�y���}w,�u�؎]V&���RH��`�e,ܝ2���^��+�8�6��� �yO���{c�33������)�x��1�\�Z�+����: ���H��I^���k�Z}�}}�0�~��,=Y<a� �JL?+y��K����*͟ldK�����y��b$ �qr��vQ�'�c��.% q���Fv>�O��'f"t�ר4V°��Y��@����>Ī�}{�����pQ����_9U��.?�~
��T�\����ÚA��}PK�X��~�yJ�d	��H�i>S���+��N����x�D��H���`su}���. y$ ���V^�
��!��2����˚��
�f[�5����m�g����Y2�>
��պI�IT��ǫ�u.�W���)�~�+��X��L����\/�/�Ozn�GNHi�͂�gg�-����PG�񒟲�^^8q�<�}3 `=���'O�	�J"�$�c�D�t��j?����y��b�S���A�[�>�=��d#�!�o6���b�z\�K�oQ;eU�����N��}�i����}���9�\(�0j�������M[̀��a�pҊ[4��ul��H����l�M,:~��������:��}�<�un}�q+�ƴ`�Z����X�|�����ݦ�MEC}Vq���9�+p�a=�B[$(SW��pk�sbmY���N�?������n?�H8��)��E��;k��O]8_��^<9.��Ҍ�=M�k:u��IK���w�W��,�,f��� I�{A��A`�M�.�1������������kl����&�M
�,��]���s^���[��v����b_�V����'��\~����%'�k*ɡ5�����`�+� ]�U��J�q����2^����1�����%ѽ�yg�Dg/U ����R�S�:��{PnK�������a���n�h_��"My��sl��^�m@�����}����,����!�L������p\�si�ޞ�N��\ez�!.���u�L��������of��F&�':_IΗOyN0�Rzٷޯ+k_�'�Z�?��/�o�.��rhp�Qi��9��®�lB[
g�(���!�'=��ȷ���_��o�nzBZ�N3�S^�Q;_^:���8>�X����W�X�F*b��nzD�m�J�L��}0���i#�+,9gw8=�u�z$��N�D�Y�c�)эX��c�e���_zl�ֻ���@�VH�4���Lڿi��v�f/� ���lI�Q���xR<�*!2�U$�����3�2�Ԁg9��]c�L4�Y͹޽�OX�������A��1��H�V���~,�Ź�x٦���5�[#P{�����5���M�7��χU;�F7�^��V����vx2��yT�����u&��c�4֕��`ךiY���8ew]�w�-�/`�ɹ+*_H��E!R~L�f��A��$�oΠ���ccig:���`^�N�L�(�F�j3q?	9�Y�}]�V�N��}���#�e(���,r��>o�~P۸;��}����	;~��zŇG�n��E�fT'�voS�A'�c�� ]�@`����6&V���c+gOD���ZD��ۂ�\9&�{"#]�o#�ĩS��ӈT�,���qI0V{��
2���0��� ��J��ؾ�ʼ�5��Q�L�dO-�Ű�����n��'�r��.R{T�O_�>�|���C;t���I?�.n�G�������/�+�Yَ�^+�@e4e����g	����v��TN���#���k�ıN��k_#��m�Լ��,,uP��-�����d4��+�`�`я�e��,Yj�Dԑ����� ��gB�|��KU"Vp��2�0�#�^�ȑE���Ҧ�V�V�;:��ֿ4���c�I���?��ߌk��[��\*ŉ�,Ļj��e{���J��&�P��dlVKq���\ީE������'��E����E.T�.��Q��@��/�M@�t"#��a7K��K��|�`�[�	x�ӶDR��05=>ػ�gG�a(_�؍�j�@j�|��1�}W�����gt��!�v�l����x��B���D��w�̡��sW�v&�:D��=g���W��,�����*r!�����].������Z��Z�����0����q=<�ё��Hq�bK����7& ����J�jh�[duo8|sF�z�w�!�
I�|z��}V��!T�gՀ�31���H�#���l��s;�M}u��c�Pe�����v����R�ُ9�0<ttY�v!8�d���8��T���я�L�7�W�JI���S��of="T�ޭ�����$ÃCwXi����|�>�c��~ ����/���R]ɸ���	�[���6B�;o��^��mo4��w2b�����g��i��'ŸӺЧ;x@��P��B��e�A����?"��|:^3��{2m�����
�؈��|t�R����?F^���[��8��1>�[��	04Ar�0Z�}9��F�\.�oøv`)}8�c�I�6@�7#@ˊ��5�^���5��?��>%h��U�;���n:o���OK~O�E:��]�g�d��WPm�xE�q֓?�t �^7}���|vZ��?��G�sy��{P�{ғ����-^��6&��ɋ0�9R�-���+4ϳ��g�q��Ă���Ư��+96���#b�ꛭ��/�������1����BP��G�WN���Fi���T�&���m�~�rW����t��	�t�D.�yNg��9�r�I���o泊�0E��d7�u�ҏW��-x��(PUL<��,�@9��T-g.%g\�-ᏗF�x�Q��O=H2��U��­�~+P��*�t���g���ā̵d�绣TD���t��v�F{�utH�N�ދ�/��X�^�M�/��Җ;*�v^����;���c�>�۬m
��s3���X��V��*hW7+q-�|�>Ҭ|~m�>�!��""���^3�o��h8�v1T򻕼��Y���0Q��v��uo��2���V�P��!'���@D��㚘�@����	�Z�����P9\�d��/"F����3
/�q�6^�A�i�(��4n�"Md�����KȜE��ԃɽ��w�������I8m����"zo��g�Z��TK��2�����H�����W��4؊�$���Ͻ��S���gt�|ˬl'_����i���y�I�i��<�MThh;��@�].� ���|oU����~��ZE8����Że.�M�L����E�ހ�L���0�~T�;��ɞͶ������,Ȳ��3�t���ffǹ^�)�ː���� ���Bn��Ja��eS����Nf����lMO��b?�����'']v�/<�?�_d��9~�W�&�A�Wk��+�,��d�pH�:I���ˌ�{���	, 9�w��1|�fu,T>����j�c�]sغ+��^8A[��O�v�V�:n��x�|���}O�3+..��υ��Տ{��'�`�'�5�P0qQ�omK�?��+)GL�\F��f,ф�^l�'���pk�H"�g��☄�ێ��>*��̌�:Ĭ��m�b����*�7��+,4�� |U|ryy�0)���Ӛ��A[�����M���.��\/�0�rA!���/��SQ�F��9�c��6�_|���CKA�Dl��Ԇq�Xg���8~2%��Z�y����f!��]���Ԍ�6iF،�%Q��a���Fx���u8�w,�~\���0���M���m��l�}�zn!����V�L�f�!Q�zř�-�LZ#���I��]�,'��nQ�}��[�Y�N�$_��'צ���!�j	)�.��Ѩ��r���i���}?�����̌��C�>κ���^��8{���V���Ë*Ëz���Ev�_^��$����*F���|ᖑc\��G�^N��m��cFC������C`�9n����_ª���T����6��w��w���׾�ة3څ'�E����9����
�Hw_���#�*}ݚ#[׻z��� ��nF��Y�2�[�F�)��){׮��Ȯ/{z����D]�?�	�Ԩ�!�m������oP&��6���jW�d�=ީf�F��4�{y�iTث[�xNL�����]_WӡJ�H�j@��"��Qi��v���~2�Z*k�c������&��n"ҫ����]уV���L��4$�^�bT���'UG�l��
mA��&�t7��p}O���q�*ˑ����H^#�ӛq�/� ���>�]"\ 9��������(��FR���&'�7��������G3���5���`?����ri��9���5a���^�Z����7y{�"��6�-�Û��z��W��IR�x�j'��'�Mlu�LeN�@���4B'�b�;A9SՍ���,�W�Lk��j�zM�|�RZ��\j`�[��v�G�����=N|�Nj�Nʼf�]����̻��x�^���:�t�]���[�8^2�e>O5ÿ�9��|D��r���:��P�Neb ����D�pL�]��Y���4j��b��[��p���n\`ݯ_���Dwa��;�5�嘜rD2�\�_��k��c��̓�Td�a����&K���2��k�!��B�/bw�u�Kx����o�+z��t� -	��P��CR�&��y��^���[�=sU|u�N���:e2�?���5�'
�f��~�w�����-��������nN,��~��G��>+h6��ѿ��=.:on��K)Y�j+O__h���	�҆"���Rn��ߏ2@��C�a���(�c�մ۬)4TZ$	׎E[D�9p�����RZߴ�0oF��n�����h<�jCѻvĸ��feɸݚ�ɔW��x�[W�)ȿ�_O���T�j	O�ZN>;�����)��O��6,�99��`/�e��G��E�a._��x+i�	��b=F�yi�5���[c����n�al�'7�K�p��[(���aC�����٭����	���EIʧm�����$N?M��FX*�t%o�w|�S"��_�0�,h�	%3W�
f 3�o�z��9�e�fybw.���/�����7��1:M�8�5���"�R�y��O>�q@�"��̝��O�^&�85K�ef4d:y���Ԥ8�OmҀ�À��~��̨a&�ˮQ�=�z��7�.P�u&�<Զ����9�*ފX{��x7m�i��������l��7.�8g�������q�z�������Q#����4lk��3p:����r���������9��;�����i\��b�����Љ���x��y�(ׯ�鐎�((�t+݈t�tw��-J���t݌tw�C�H�{�9�����{\k\�r����{_�8�[��bg�k�T�8:3�>�qT� �IlU�+6�@f����@��S��mkĚ����U�|)cU��F�ͫ8�X`�sEO�OV�̤�J�<ƹu`ۘ��K=��
x�}�){v7t�v� ^D����rC�v�Ƌ���<C�?/89b!ٌ�n��F�|Ϟ�g�� Px粀��KĒ�^{4�����2_ch9,�v�����rO�5��-�NN{Bk\5R�dQ��D��'NW�1�/[j�k�}(dͭ�jCG�		��4z��d:	��ž�$r�5���5����B�YW��@G4��kTD�'�S1�!~�/� 1,rlO;ک��J���M��>2�&�\�m/�^�����O\�`�s��B����$̿����æz����HD� ��K�L�͆��*�H\����lJJ�����nuL��\���'o�8�@֐y��Y�L4y��qa��p���ءYQT���l�y�����*�e����0�F���K��[W;�=c�V�xh3�oK���LOYp�p]��>#�Mד�*���	�mI^���l�e��֢��msx�����`�P����,��AS!̓��2w{J�E-�#N���(S��-���E'�P-\3Hvܩ�׬��)��: ʈ2�l�`����j����!av̳-�X=J}���+�~f|r>�kc��`xYl�C���В���P!���g�uA-c�h���6�}���F���ظ�����W|~�����ī�*��Ric�SA�ϱ�*����e�s���P�x�yx�Ax���ڗ�W)�L$iQ�0�����S���^����K��T�7\���vi�D�ު���,f���+j�����w�R{C܇����0��b	[<c�t[T:ۘ�4fSn'�O���b��b�Y��\^�ɽ7�,�R	���ӘT}+\�ꓫ�U�vB��qMX�aXE��m1�4��ʢ����Q��A��
��wj�7����<1;�B�#y>mY����@}�`@�]��#�8��]y��h����`��힃���K�-��b�}��W?mg@�!������;�n'�a�w'WQ�@�k��ƯD�����,"�mV�t+-J�W�"PhK^��4��z��=��f�������g�dH��>5W��Ş@���X `1&�$���q?&�?=.�n�+ޞ�;y#�v^�R�/̉I�fkг�aY_�"��yW�d�Z'�N1�����P=��<*��w]����z�ft���>�g�� E��׻��];�r�\����ٺ��\�ew��h��>���Z��]�{��̸�BO�M������w��cc���qי�u�olS��mS�}t�|s�;�|�$;ۂ#��iu����7_ '0��ADh�>�Pޠm��GK"n9���x���F���Y�{��e��ʥ�0%9��E��O��o�x����L6[N=�*؞j�$��Dc�9O�^���	;�L�T7J��o�3z����;9���պ��a�iႥ0i��%E��ԟv���!}�6a���`���;JG.9�u�(ؼK�fT&���M��r�[岺�8+��g��,��L�b�}D^�O��DT�yHB�%3����,�mk�ė�#�U<s-,%��&�@�˪{Q��R@�{䍶�����VՒ�{Y�Ĩ�RYU�<F1�}0x7.l�R�7�h,�J��-9����7��Q���u�7>�c���h��[����lRe�)�_�/G"�
k\V�Xʣ"�X&�C�<��<=��oXJ���=����A������n���ò��{��0�4p����w���������@s#��F `ۋ�\�K�2�����Ը�iy\��̒��~�`o'P��g"�ݱ��BO�7�L�w@����2ښ�X��������vKW��e���c����<���5T]���`㠯��u��ᮊ,qf�"�v+�����b"����U�'��1��(�:O5.���_��5�r�������-~u��� U�lqũ���7߲s���$��ޟA�ds�(Y	�I��W�v�D�XE滈�+����w�%�7wH��g|i��ɧ~�y�1 }e����;��4یǅYEj'�;H�-S�A�r�\z�*� UvT�-J�|V�k�p�6�;�v-]�Ƴ\��8�$��Ў�
8��n�t�Aoz��|�׫���0o7�����Ԍu�Q ���]��q*�Vּ���ʥvp[�d���_���a����'�NcS�]A�N�--\�zܭ��a|ȇh68�@��e�Põ��n֯����r<���! �il�����U�2kû�k�%<g��G1ݴ��V�ˡ̣��c���M����u�`5��YjQZ����_N��OQ�D�(.�ww�c�[����ى��@�U����ϧ��j����5�z���5}}x�ko?������,�C��҈����<EG�כ1��#p��8��r����ǔ�ĝ%�6<o�ÿ6���M{�p�&��;�c���N�5��v2&Rn��T�ˮA�y%�X��3s�9⮖�˄���x��Еm���%�b@e��]1�������6k��
���tO_� ��'(���"u}c@�E;UH�-�+�U"�#AYq���p׮<dڦ�n�3`	i�3W��ç>{[줳�c�J�Fʥz5����� m�-$�i¿1���h�D-@�兘�V�\�O�?��D��#,����&�'P��V��b��X��|�}�ml{%|�&[\~Z��>�gy&�M=�Ԑ8*i�ZM�݊���4Ot�ӌ�3?�VM1J j6]ɽ�s�:3[)�w�.f�B��ڷ�v����\|�]&ym-��ꀩ���#KT�a��RT쵔�^����gܼmm���^b�:������������<%9�O�ا8�M�GKSZ����m�Թ�i.�T�}��RTT��K��I�(�NN�8�7 U+��N��~�-��ߜ���yp��]�t����r!��Y�Ō�����(�"k����ԃ��V��:�A��{,`�-�<7��\j�y�~P�}��Ǭ��*z�c?la��x*��M�����C&��ب�sT-QLp�2~	�ѱU����'\>-��Z���x=e'>b�������"P|<(�>چ髎B�F-�Jˬ�� 3��萫s�8#�_�,�������'_��me՛��m���������;EJi��ȴ�bG��iYD�^�p1���׉ϐ��`3�l�}IԩLTӦ����T5�e}ә;Q��鷚���ft�6g�ר*ʏ���4=�gY�s�UU]%��5C~� �Y�~����O^�qOx�ڨ�w���T�`�K�R��+mB��>E���	r��g��5.�[,���睧B����;���n^�~7��ad�@�T�Mq���/��O��Z����}�gs��~6�4����у�/��Ca5|��T\2�.U���g�?߶��o{v;�`�e���)f�-��?*'>�/RBc������$�\�K/�MX�Q!�WI��ސ�X~�gO�P�cZ&z�H�e��&<�nr
z]̘S}��ቹ�@�_ER��OE�B_!��)S�31>��V��n�`Q�����h�J ��r�� #���妷�������;��g���
^�!�nPн^���rE�2oj.�t'a��+n�s�D&�n����ߋ���*��d;�i~�$8�{�d�!up=ggLVsRPH�-�k�����w�w)����u���8�0 �tT<C��N�rI�� B�J�~���#���h���PK�#��5I��������!��Y�ߪjlK^�j8 ��q%aD��7�zST�,�:g^e�[q�<w����<�0���At��2��x���#N4
~�cr��3�A�J���ױ��|^0�!�<����˃��DGB��X�o�cY�x���/���ŹXQ�x-�����:����Ad��?�����\���y���l����-i_�!��I�q�n�T�7�5<�Ĉ�C�i�t���ܞ7���os���$8�������}T�������noKXΡ�}5�FP�ƣ<�Ӡ�?�?
��:\�q �>3���XΖ &���ڛH�zĭ��n���+UQ��5�@Dp�����W�J�~�x/q�?����7hF�Q�X\��R6�����ՙ7� ���f2=0����v�b��C7�ݑn��N7������:BO��7�;����⊹�&��w\t�Mrk�n�;�v[o�^}^=�_�D�>W�<k�P9�K�	tr"��}�Me�b璵��%�l��!�<��oϻ�T�	9��Y:���r�2���0�H �|1����7��J$�nC����7�;�i2�=��b`9�|���,�oe)k�-�ᐑu�\��/M	���v��j�42d��;m�%54- &%Iׂ�����gc��ǝb�H)%��4���7O#%�r���b�� ٕgՌ�i�a�p��C�R��A��V��t� �1[�ӯq(� ϟ}����i�	�S�+�JZ�!�L�F}�ڮ�����~�-��C%����+r�=�8(�bk���c�2/�Y�au�9ߔǬ�5j��
�dծ$؟�g	���55B������/a��V���2�&�Z�z���j�T��a 2�S�O��:�]�	Ӊ�"��"�1*R�"���enۻ�0�C/;Z��`sP�nG�iаAK���՘�� tK��j��oٴ�;+�\��w�^�Դ	CǄ*�!��ñ��:��~kA�g>'[C�'u
�Զ%�� k=WmG��[P�5s�W�+-��Qn���Y� +���#\����Ep���w_�`�/��ސ^¾�6��H�m�� ��k�SK�?�kvVмY�j
�,FH�
}���a����@#$�8G��ЀA{>+W1�._��r~�2�՚3N���f���5[�ڧ��g����k .��}p���+k�l*痆v�+�����io�î�I��G�˻��i���6\�2O�AE�X��a�{O.�![�A^*��uxU�rQ�ǝ�4���4�Qq8�9���:	������G�' h'��)���Uꇠ��C��֛B�l�j�M��.��@�uF͘���z�_��Omך�\ow��|lG������ș \�haq1�{�~Ko��,_lf�3�{V�3��/gl���H����'Ь�[Ue���D���3<fo܏�7�x�ʩS�������Z��ԯ�՛�W�6d&���{���ߊa�4�77z�T���z2_�z���׭s��@��x�>$Tm;?�7�d�͕?mce�k�Xp]5�e�CM�s/�\�x�f��,�8���4��)IPSQ�,n��K�>��p� �=�j1������ᜒC��(3&����zE�A�:�]��Ԭ3޿*�*�6Ϩn@^)ހ%.�9[TxՠYX�i���iq�+E���9�7RM{	�����A�7�v{Z���O�����6b@�G����t��R��rhc��մ+���r�tZ�ߩ��=���Dy��=����js
>�g���F�qHB2�@��e���J=�.�ϟ������w22�9U*����T��@��O���E66�؎�k���M۳����kt~���Fb�j'���%�j����M9�?+D�����:<U��_۬�r扳���E�OGl}�C�m	�s=tf��8	r1U'g�R@N��N��V����oh�����w�AB�r�䐇�rsrƢY77]��5�-�O��D�_��� ˇEQcE:�3e�t�D=�G����,�f,c񶮈��x�l��h�u��l5H����4*l/Zl�!�����#G��<95�茊f�HC<���r������Q����)x��ةb�Zַ�VQkë�b�@��<�9+'�}�E�3�!���f*O���i%�����j�A{�j*��"�y�ۛ�#�K�"RĂ'�Y��o�dL�9�OE@ou�XD����ղ�^�������A�	HW�1 ̏���iU����
Ě�E�'!!$�vf�O���G�AY�pL3߂�S�:�_��s�$�މ����ݴ�!�������%<�����d"@Ԥ�D	a��� �@e�f�t�U���,�(���1u�2-��8}��+��C��Z�7��R@�#/���<�+]H?�j�u�t]D�%fA+��XE���V�G▌}Db��y�b�����w�=0FUQ��-���y �|<'/�ǔm��"�K�޺���}1]��&�}θ��`�r��bJ$OZ!�-/eEm)C�B��K�j�,~�'*ja��5���T��p]�s��܅0�]
qꓬ	���� �h��ѩ���Sl�c��y�Z�C8��v�Џ��(t>X��re�5��i���D�~�Bԝ��0��_׭��C�;��*m�	&�^�V�޿�{g���`�x��-|Q�ѱ4�&�y5�X�P��}{|K^��~������v���,�d��gkV�ݝ�*)-7g4~4*o�3ԧ��a�gJ��,G���!���'�Ip�q�} �WJd�Q��1��jy��~Mb���.-�)9֏�Tξ��j�i�[�4���]��[N˟��W7$��d��؅u�ľ�ޜ����3���^!����K;��$ �_cv=za���xW��u�$��y������w���ƅ�Ծ�k�M1h��Y�lM�� mv��;Z��J ߐS���%0 ��-1ɰ�����"�)[���?j%�`Ҹ��GY�^k.7P���k������V_t�a~^����1��;��Q_�l��9�|�@���f�v!���l�Jv8�J'~BM��d6*'���(���¹�i$!V?�U=�Wj����f��N��W����6M0q	���M͇���Y(6r����'T�m����!w��[�g��Z	����]p���5��e�8����c1V2�I�ZL_�=]�e�nZm���x~�s	��`�4K�	Pi3�z���<�8}��#��ėk������J�~��f�h���ҷO^����R{��^ON����p��D�8�N�g�����uң�����Ga�s�6.�`��a���>�B��_�_>����C�����_��s��=����9���?���m���m	��Ĵ���x��S��������m��~���"N�o�*�{�ۄ���+
tZn�W8%�Av$�%�"��S�?�_*Zȹ*�|����70����m����0���9Zdv�t2�l��l����1J�\S%��ReP'��R�Z� �5T)ʑ���n�����j>��%���-�*e^%��k�����^'��uV31�j��%��:�l��epVF�J�WhI`��l�ʕ:�n���棅�r�O�?�_n�M�z?��m�?p�c�z@�*�,Ƃ�5�F�Zk[ܜ:�\�[��T����ؼuX����{��E?��^������f��N�Ŕ���=�-t��۷��9{��H;�#�b:j)��587����௦���q�U����!����w]��Y$?�п��`�%<�%�<�8S�;�6�{�wfց�Y\{Œ�H�V ��e��2r)�b���_tA�r�Fu�(3���P�sӅ�D��V̈Q)�&��{O�x�].�8��%�%9;8>�9�������9���n~x-��#V�T�1���;��.e�n�x�r�l����%�B}�r�%[_[+,K��� ��������<�O�%����;����]���{��	ܵ��k�l?j�I�	�kʪo�v�w�7��F;�U���������v_�;I���)`��Vs^���T����1?�i�-�@����1��֣<&jZ���"�e����(�,���-�ǏF��n��W�5�LD1�h(��߻�Ф��@�d�����3����?�g��ٖ��0>�HgX�^)�y����8Ѐ����-�[�QK]��>�3�J�r手x��6cN�:Y���V_,F�I�6ş7��O�5.��N�-7������aڃ3tB,��#�r�k�����)��HP~7-��<��aCRjn���w��=���Sq<�7��|F�C�y���0 v�J�ڤ���>Vȩ��5]D���	w~x��?u�?�%3��������ѽTe�A�y
����Q~W�B>�g�k8bD�$q���WOmd���>�9LJQQ��4D�t��zg"l|Ϟ�������Ab���M>�>m�����{��4�xu%O�*����'�7'N�WEA'1,D�G�rKڈNOxo��h�*�3�����3J���*����%��t�r�ֳv�$��f�+3��s�n&f���<��P�h�m뤸���ׄ��/�S���.�`����s?���D�WN5�1p����6=A�YB��ůq3ދ���P��s1�f<~E[w���^/�L\ܲ����2ܻv)$e~���D��=��^*F�L�e�eEn�\Ϗ���3�H��C�qY�e�U�ɹ�`��60�y8*T���q�r��4��/^�H�]��Xd6'��vO�p��X*�������s�v�V�4�jM��i:�n�ɟ H�qb{8���x�I���ˢ�`	K&-F��>�W���s�������O�3k���vRE/P�ˆ��&���oAd��ڮ�=�X�$�@�zV��ћ�C#�Q���W�6SӅ��}��+:�4M�ӫ.���i�_H�[�����M�^�����^#����Z�c�s��� "c�l�ĄF�yÆ
�AIJ�ȿ� �ޠ����Jz��O>�;�W�D!�@m�Ʀ��O��k8ōA� :R��8G�v�'|1������q�����o˿G1�@<�8��u�ι��#�&@R�{�L����\枰�������^=�N�-	
�Z�S撇��9������ge����њ�-�� ~��ZDQ���U�Ga��P�𯱁������"K�Y�0-P����������a�e\|�N���\�K�����!���\|"G�jla��C��Ē��Vʨ��<.0*Rn���al(z���/Qi���[q��6D��#�v���/�Ζ�P�i=�� t�ä��r�u̔=������<�V�}����\T����j�^�<�eE��~�����.}��U�Y��`Y��$�����`�m��2������p�������zk��|�JN��?���3o�K�����Ukv���!ު����
T�k�6�f�f~Uˇ �
$L��N{	9<=�{�iT+��hkJ/#W�/6��3E�~���a,#��?17�=�e���i��f�B�<`rc�Z������;�{�:�}���q���^�Z�p�us���
�}>�����6��.� V �}e'���^���^���(ĵ\�K�o?0���QJ�"'R�Ө�C���j2F�S�~��/�g�7n�6l�Du���&[�XLNF�oDx����7�2�����>99e�@m����|��'.y��rt\Ty����쨭�J��iz�k�%���͹]f��T@����\\ܩ�7ݫK��]�����R?�+Oܟ_04�l��1��!�hwV�wn/�ht'��Z���o��(����?����2�g%UM�m�T�xL1�Gq��|�aBB*��χ�~��j�qJ�0���o�����#��n�g�Ph(�&i���4�\,��y<����6p6Zz*m�>y0�L64��(�(?�Ց1?���h�܂8�M,L-e~��jSߵ��2MgD�gK?��汦4�ġV�U���+���?4��u�3��D4�68�X]f�������Y��8da����G~� e��T��0Ik,���U���V�����s�2�SdÄ���os%��ˁ����ja��l��.����vR���0l�a��ǀMG�oM�o�
��T��=�w�����?���/�6�kCڛ(�Y����+ə��_m��Y]í�o"�R���S���8L$�K��1�g
�Ǝ��cO�,��W�'2PЫ.�u֤ok���b��� 9MOcI�����;�G2kG��nθޞ�t+��^��3i`��5�0�G�#���NGޅ��J�K�b{�݈U����_n�]_W9�:!����H:r��LK�xF*&.�Z��b���N��9�k�eN= �����ݟ�&���o)��\��o�����_��e�^!�E�'Ý��4 ���ZU�DV��ư4nh���L0o�$����r8��%*�D�䦗jTu��h�k���;�;�͵�Z����4:���ׁ���.����0ML�)��M�'`{���Q�<����8�����H};d�#[�JKlj�E�_��G�S`YM�����9:�5��y�e=O%�%7*���_��>�$�u _�&w������inPmu%sp�ܚ����h����	ٿ�-�L�,��
�.�v,���ڣ$�0�*E��>#p�]�� �a�Ԏr�J��a�Fxk:��u�}q�~��S������>���@�����ܚv(�٨<�q�:TV�aB־�|>1si�w$K�[p�_��l隸&���;���@V�zL��pO��wy����������av�Q��
ǘ���,�^э���Y��_�#��"��j/��쾼s���3�	�?:�9��[�r�t�J#�3a�;�; A
�{S��qP���'cP��ɦ���)�%w�=?��I�1dFŐ]�͹-�h%��� ��ٶp�y�34`�T����*8W"]#r9���a�3�~N3F�3��a�4�8����К�X��J�<���h�4�ح�;(2f�����Xoo��',1�1��R���`pO6oh�΂��{���x���8������|��+��H��ս{Zi��!�F�F��|�
�H$q6�{q"�*�]rx�x��"?s�Ɇ=�0�A���D˺��!\tSx��mM5"��U����:/�T�ی|�b�f��~I��(��[�=7�a�fuxpd����`%wadI�~���/(]� �}�}��&�s��r/[�,�������PxJ�ׁǂI:���C�_�3��z��B��=�A��䯅��8��ҩ��U�8���m�����=���HZQ�[�n�J��7���	����C>�D�d0�)���n�g=�`H��M��Q�د� �GC#� ���-�Ă�cZ��~�_a��/���E�(�d��G˖dlPE�^5�ly$�e�u3lv2��>b�6G��M1ٙ���̞��Z�-���.�$Թ�E�~>�����[m;i`br& ��?�A1��?�#��e��K㸃�~��/Wp���b+Yp?�L��0L��|A���nr>�Oa�Y�6��<� ��������=��K�{ë�N�C��0���̉�E�|t�5p����Ѿ��q�'�-���Zg��f>���+�1��8.����T��J�z��\���oMu� Gz�i%�=1�+�N�L�X�%Ϳ	3�6^���� jO7#����Ǯ`�76�ے:U������1@����7��Y[��K��aJf;n89�[+i�*���:�͗c��o$G���f�4U�@6��� Py��k���#S����5�o��C
Nr�'m���o�G�����#B���%�,@�'��`�;��M	h��:tl��&����8�p����r�7��7�%�e���ذ�Gw��`�M��Y�9H��G0��Fx�q�1��4x@c�U���ש���#ѕv)�4��3�_�N� �i�7���əUNw� h����5��c�}d�B�����7��^Y�ا���4zd����ʂ��W�;[!�"*M:���N�M6��xX��1�9v�����Jq�WȒg3�ް�`Y��ĉq�w2��^�/_�ݲ�k��
X��)�չ�Q��tU�N�צ��9��c[���W��t&�:� ��&��r�3�_����}�˟���]Xk�o;=;S�AeH{�JU-�����W�%l� ���yk��Q�ewg@o$�kSa�@s�>/�[��Č�>�W-�Y�[���=��M�:ّ)�	,��- �1v���AJ�����
' �Ï]78q��hc��8
Ց�L:C��6�[x������r�Hpv�'n�釈U�W�k��+�=�:9t|	TZA�A��w�����0���s�ݥ�I8Ư��p��M@�&�a=�Nٛz6>@��#k*[M�mt�D�(Y\V]�G�w��܌h6W���j�	M^�5����f�
ʥ���#�^�#}��`C}��|'AQ�R�`/ѽY���U��k^M)`r.�6����Ɗ��x��"�su��/r(�7Ԗ[U�jrࣱ.�Nd��S�)����[>J!Ϗ|16�b�2g�C���|����.{w��V�ZZm}��f��VQ��#�r�)���������N�+�T�.�{-�`������@�G`v��\+hK����{�l�)֊zl�pɮu��f�ź꿩�	���	�V4��.�oZ��6�|a����O��������ߘ �c�7j�+��Y��TDrEB���J��k&�E�P	-�s�ꇄKq���7ONT�b?Q&:�?5u�=��?σ|�L�+(�}k�KC&��^?i������>��I�bB�������w-O�[�m	B=4⥥ۥ��wN���z���;BX�X�G�������-31j���j�<�}��8~�&�ǿ�<{�9��:�e�kH��$�8��/�H�q��W��X�����nn[ē�m��Y�2�>���HRC�������{{�Q�=��eB����לQ/�y�(�x���R�C��#�Ta�ɴ�G�ܬ��$�ώ���h\����4d����1Z�&u�ĝx�<<鷐��b���8`�W���)�x���w;�G����f��}��F&a<�+`]e{��Jnj&��@����!C�ڐz|w$�NF��]ԝ@�����Y#> 7޷��<�p���a�,�~y���%e�0��;��	�Th| ������2Z��pz?y����t���O������v�<��Hh�X�����ݭ+@H���^�M�,Q��/�.Ql�!����`�p7t��9B�d�h.U��Y5M�}4݈J�Sa4�|�ws��Σ�}�קv��Z԰��O8qXdM�>�#������}��H\�W�]�.U�BD���|�kSMD/�����.6v�+8>�z��Ԣ}$p��,��H�)�5�����ɔ}�J^,�S�����+7���&�}��#�����vw�>�m�뛵�S����� ��]&�d�b �̈́>1������&Pc�_yY�Н�;/�L��Vְ�M�v���eT�#��O?e��T�$B�-�Sv���V��?�Y1?��	f���}��ڈϰH�SO�����)J�#3?�@�@k�{n��wd,�D�Fc2� ىHdN㭯����&�<��\u�x��\G����H�V.�>��13;��z&=��R�������nW��EL_؈�
�1(v�W�Y��] ����(tQ��@â�7�Z|b7^[�za�3� �������7�k�� �ZŬ_��
1*v]�P�-E~A(ބcܐ�&�M�8�b3�l��v��nf�q��"W��
	�oO->�\���*X�A%~�KY��i6!����_����"�F�"/2�6!i,��W��z-3g nŬ�;?�Z��c�Me��
P��fH��GU���w �JG?�T�F�ĥ�Z�2�8�}]ơ���ń���^j�h��ED��Qo�qQ�H�v�_������G��CvB��IN��8�4��~%�e_(�?v���ul��9�Z�R>�����U5 ����1]J��mmf�N�!8ЯZ`�L��?C��h���RU,XB�\z�.�_]�=a�jjd�C�� �� ��|r|����fmi����jq�����5?o�IQ�&O��եp�%o<������#>��w����! f�F�@���*��C�h��))�h��Po���5-�złb�g�3E�v�k�%���E����8�'�JqһCD����[�KV�b���.�o ��*,�*ވ�5�������������jU~	����~��!G�e�� i���~��|bFA��G��>P�6iTyx_�-G�R�[�e,d���<��>�ְ�����6n}a.��8㝗�_E_�l���nـ�`����^��;V~_��X��z���E�I��		�缄�O�Ֆ�~6�
��M�3��(w�@�m��|F a���1�
��qh���?�J;�>�߳��{��rodi4��
N�$���vA"��0Ҩ+�*gvNq�NO����]m:��F+� �=���U)���� ��d�D�
��@����aNsD��x��k&�݋u��5�������W�
DӥGCHElq�<1��X<5W�:W�O���YmyF'��n�q8!^)x��Zy���+���8׋��tƍ�K�V#�흾j�uͿ�V����{���s3���L����4���[��^ܐJ�K�#�}�G��O�` �\J|�x�9���̱����h���|)�h�����'/��}�D?b<B���Xɯ�>��!�	���K�|�t� 9����%��A{�d�
{��bGc��֖nX��n�Nf��/A��=�k�T�w�Y^��*!�~�޻N#!��U��<a�i������w J�sө�'׌��{�����s�w�7�F���)��s�x�T>9y��1nD�̀=~��p��~�э�cf^ޏ�M�I�_��T�{DY��sp} q8�0BJ)s;�(��T6]�]���.2�S��0֓�cp��3f"���a�	�_�@�[�V��o���P��"� �X���ʛKS��![���"兪A���~��ػx���[T@�j.!4}|׊h��d�'K0J�W���YHa�x<ZM�e���`�x7? ���5E���ە�V��(M,��?˴L��;ֈ�y��4HÀ�N���<�G^�
��t�r�&�݀<���r�E�YE�W�VL|��N�q�=^�1s����x�e펒m�V?Q9�7�>��#����.�C`��W�k ��r�H�5,����ry�*� �{��מ�2��C��x583�m`D�_�i��7�K���X��Y���)�SC�3�=����@�o��+ӈ��O�"�N����?~��`Fs}7��C\��b��Ԭ����7Dn�r�H��ĥ������*�A���|E���&Z{sp�hX�a"���^� a�境M|�@ք��<��qH���J�(�F�/R��|��۩Vfe����!m��͐+�	IPsrI�/A������i<�Y,qӫ�|���i�C"7�� B� �Z@�im)����� B��Z51A@sL%�#�и��Z�F����O�G�	�~a�
�(zf��1"o��(�t>l���;<A�w��r�����ƾϝ�V�x�w��P�헏�bd���=�X�釿�!����B���#���)O>������~���Y �L����X�|�g��m�M�Iq�t��J|ш[�%܂�-黶ϕ�9I�8B�qB�J�� z�"����s���Ad�)W�f���`�\�|�S�R�vJp�����hBba-�%���3F�3�q����/��y�Ǟ`u����I�>u��͈���Iq_YE�{3�N�	2/����(��,����oy[
��h5,.��̓��"|ܽ<���\�Ѣ��.����Nz�U��]��n���[e�$��|�K�k9p�ؓ�d�d���,&�O���*ōs�&��!W�Vαﾛ���4k%����8�>�~1��L�d�e�"�x)f]Gr�*��\x���U����5C�F]��a�(���ۿ�ڛ�K'7��1����J.M��Z66{o�Y{���+?=5�ַ`�`�<q�=91|N�^ C�>��г��v�9���'z�Y �8���rD��*`!��󐅁��~�2"Ÿ�̢F�#�����Hb#�,�N��ϗ �w�_��辞��&�����"�`�S[��l��è3�Wݣ1��RIČ\�QьΡ��d�O45z���n$g=����8iPa����FEK�=2��1�A��@ęm��GE�*S��uw�X��J����֩a�����B�B�x��Pr���Z��%�i%:�Z�^��y���+���wzE����+�q�	��{R�������^ ��;�ڧ
_j�ڊ�sʿ�TX�Y��TO��8yu��@R7#j��:�Q�Sd�`"��y��{{|;����I,q/��V?������'�?�UR��a��s�^Y�����-^Xˢ��7�/7+B�'�=��dt�nG��.����<�Cz��8�R2hd�M�5A����y1��.����� ��,t �(��}��l||gs	�?̨��<�7}����{DYj0K2��mM��5�5SV1�2�e0����Ce�G���JtVUJ�|�WG]�I�=X��Ś`�W@e�=�?�����������^��~�hԉ|V`�FwU�PD>�~��+ə��UZ�����[:@t�T�ao�I��Lt�#y��æàk�!��n�IQ�o �ʔ��ۧ��d7�PV4ގ�
���L&���;�ec��#p<�����`�k��@CkpZy�{�m�z�.wҌ/�d�������!g����� [�_�u㩏�q�:1��|ޓ��Q�m�JN�Q�k��z����x���v  _a� ՙGTg�?��f/��S��ZW��X�j��-��,-5λl`{��C�,W�}d�{���#%+�i|"�� �PJ�\Ӡ���N�a��!�:nǇ��?2�2*��i�@��w	��!���%���.	��	��ep���.����=���{��Ś�<�O�]�]]�qb��B�|v�.k�N��F�R��s~&�K'#K��\�5��_�4�=��G�h`u������S�v:c�P��3z�JYa5����'��^�Dv*�Gŉ��Y�Krn�b������-�� ���r��^;C;�'яL�0rI��;�&�%�A��=?�������؋=�Qy��:�!��bB��G\1����"�w ���?��ňW�~�F)���W����t��x�+B��%����k�푨�5�J8��tr�'OG��ۓ�Oہ1���b>��]��q���կ�Fw?oG �o��{��.xc�ق�[A*�⍮8z�1M/�����Ϭx�O�_Hɲ~��O$����ڦ����r��6Ѩ�� ����cҒ�~{����p#�㧆v(cSPd�ǌ�����
�tZ�q�l�bDO�_���X����|�`/�,o�J��=�����4��0����g�N$`˂�o;Qld�{�j��b��:����I޹��������_A;P_����%8~$^8ݬ��M�]"X�У�t>����ن��"y1j�v�2���X_=�3#B�1m�}���f����o�_��ABq�Gr�Mpe6,��=ڰw�L~�p�u����eb/%�����ވ�bbh�׭��<�'o�A4@\2Å�O����4��Y����
�|�t/	�y� q����=����^���.ys'ZD>܄ܯ�7~��P`I� 5z^s!�߼3�J�`�浢)}닍L�Re��8*�UO�t����:�}�f��N�k���p�#���M	 ���:��l�c�;��%t��F��:ɘ�����o0��:�ݹ�'���]�zZy_���^��Ν��mS���4��*��؛��,G��O�-�4�0������j�!���-iH��q��6@�9���X}��rx^-��zT 5�&J�y����8An�u�@t��(>�[�-��#`�ja�!ʅV#��:#�!0t���n�oPH3���n%�����d�y���ۧ��O~�U;�M.��R_-k���)�⓯8�[���[�/"��ޣΞ�T}�dLG������%�c�<u��F[���b��j�������ܲK<�қs���{��Ҵ25�da�ch��#-ӣۃ�kq��G����5�o|FK��_�Y�yK�:I��i�� Z|�������K��S��u�> �	��P���8���ő@Y���x���v�d�����&-�'�󃀇sC���ذ�{��ј���V=>׆���P���B�Ųa��~��}&U�Xo�7��]t84{]�Ǒ ��;�*��5@x��udv���y�)�Ef� bꦵ��78��G�?�,.�G��`l��r�p�3����'�"�!Y�U�7?8�sC5��� �5k^ntF���<5pA�-�_w�^,�b{'���W	ᄶ ���޺���7õ�YVyX)aK"��PҞ}i����b�����3)������xG3t�����)�9;���h"���Ҧ#r��D��u���ۗ��my������%
���S� �C�p,�U�)���1t�)������w�Lfy�T��ǯ��G:�9;��˾����|�q�ޓ��(�`�_L�?�&W�Q?ȋ������K���#�c�����#���#�g
ۏ�:��ऽ'�w�+ݡ�+T���uJ�a��8�3B;y(���Oݍ�u��/��P�7�j�O'���WTG�kFݲ�♐-�¢�ߞ�����ɒ���j��Jɍ�ƧY>��^4~�V�d����e��^G�Y�����fjN��'�zNΕ����� X"�%^7Tt��R��wZx�s��;g{��f�Ӟ ��yr74��x�=�Y�����e�ޖ���Vk�� �=�@�������Fpf%"r���r�>�aT.��FBV��:$�I
6�h����aN�Ym��r�/�s�U�4�7���`��(˔�UULº�^`�6�cm#brO��|��PX�!3���5�ƅ�3pʂ�Ü4��/�8=oM?
y��r&�^����Z��(DWXm��/��\�;���k������dh�y�K?-L�#?1?20,
arΏ\�''���ޮ\7:����gg.c�E>���x�@��芀y��0_�v�g6����ZpV�ۢ��:���3�7j�O�����$�UMMNOF�_�v��"� @|	wgJމa�b��"[_|��%��ro��o�j�A�I��3�ve��E�+x0%�=I��A��Q]{;�ҧ��/�wK'��H��`�>%����c��QQ0T�c>5�4机��S���~�B�]1h��o{���_<��j�K3�.��0/I�j�
O���I�u�D�ڗ#�F�!A�7Х/w���#z��
��I�yS|���+�]k�5�~�0Io��D�Rd��y,h�Mr9 ����Մ�@ˍ�7�_s>���k䝵�<c�sN|��I�?HtD�[�@Hl衋%,/��v����x�n�`ѕ�%xV�CWձ�D.1�PQ��z/�ݽ����M?!�?��-��pf!w�}#�·s�vs�l���͸��ˇо���9Z^Q#�y�r��(cHH������c#@��>L).��X�e�X)O��P��6ƈ�
ٹ�o��nD��&���?�D���׿�`��H�����w&[� ��v�i6߳a32	#��z��4��"?\05#_q�N��	��;Rh�ư�A���n烒p��]t��$��R�����d��Xn��]�(�%O��
;�B�^�T�(��aދ��y�}����	����"��SEu�,z3���ac�������fM$4r��9�y��8�����V<Ui��4�����9϶�9��Δ��3��u�v�J�<���l��U��Ϣ����Ri����8l�Y*e�]��W\�۬�YV���^�Q$ q= 1T[\RIFô[��Qd��.]�.��E1���S�ƷS��	����	����܅c-BC=���-�~�b�lD���0���b�Wt�L�� M��
�F]��OtX���&�}�V���a�W��ƫ98��o7$��.���:��Єt��7�����9ݼ�����gϥ��;m��@�lLiߣ �=�~�� ��	�
�]�D��W~�+)B@���}|���w��Sɑ�֫%��*֞d���T�ꊵN��m#兹�i !3jQ)�`d�rqs�s|�9X�h.�V�0�3Z�]<�xő�:08�F�.��Ay�Nmf�����
���%�K�M4}��:����!/�3c�b��F�"܏��{I̋.c�M�t�ʗ�\�g�g�ӻZ�!yCKF)gs��J�&^��:Wٟ���ۤ����H8��3
ݤ�nķ.�U����c$ꠣ�q�`�i�A-U��"��
;��v�ӧFC� ��_���zs
� yԑw�Wi7s�3vp��v�jN�x!�#���V@��ǹ�/��\�6g{�����v�׀��"�����f�"���н
�-�+ &��xB|MG-_:�KF�b��q��P��%o:��%��j����?w�Q Y�̻`�f�p�Dd��tO��C���^n�m��@�h�+��C!����}��<��q����JBn�7�ڔ��)��m�~>���3&P�u��p*�92n;V���5š~����"�����ԍE.E_�ĝ��_��k�����r�*�^�X�����81���}@�vP�����K�����qqnp<�� �_�QUe�o�@N27,-T��F
y��;��\+9U�nb"1�QԦ��,����e��d����8D�Y��HXO�j�1�bo܆�j�Zٕ��8�H�|�Hd�b7�Otj����U��F��x��ſ�Jq�V@��iݢ�:}���T"�����58�\5�HM,�I�@�{隍]�5���v�sl��?�N�㯣�d&���3��c�g><���M�$��3�8�'!���8}�xK1��5��-u�}�z�����9P�<Ӄ[�_q�҂�N{�I�'�U4[�Ot��7Jy�,G�����������
9@1~.	Z,����g9ThP'[T��U�`���PUݙ$z'�)�2A�(~�WS�z�o�gFe������A�n�+�&:&�{h��8�70�W�`?x\h�<&�Xt$}���y�Ͷ��BB2E�Kv����\��h�O��A�sL��#"Ũ�[,���]���9m����|pk��Q\�98��Y�Sc����/��a�������'�@�H���W��������G7@�b���YLM�{D ��0F��J|���m���@baQx0}�x�R^ L��7/�,���1�ja�2
���z���'�2�f�)�^��ts^ʈ����[�|�Z`�+�K�$�f��8pp��]��S/��wD+�Ӫ���)�x���Ʌ��*?���R�6h$��I�k_�Xl@��p� �vH���靽�GK�.����yȩ ����_�AY¬�z��	P`-Ԩ����`����چ?�_jR��Q��RwK� Ȗ<yp��nT�k�y�O���[��7Mo�9�t�Y܎�ڎd�8Ȑn"=��S��o��ڡ�2�ꓳ`Ե1��B܀����Y�������9��g��;����@C"w�!$����*�7P@'�� ��6�2�����
X���󷓮���vZ����8q�������P�<�P�I"�L������H�[�p��7�(+7G7�~^�����R��Q���<T��H�po�//W6|�"��4{8	\.N�'�^7~�>dT;��U`/���ỉ���ͬW���K�t�n��w��5��x;~Ǹ�a?��@��7�N�D��J�[^�u1
��EW���e)�i�e:쉻�8�0���w���M�p�ć��@��@o:%Es���U�ki:U��"ܖ^QM8kgoV2�C(��9�OS0�dA`�a�elz��΄�֫]��/3�	6�*b��%�,Oæ���%Av�Zk����U6���,���K�RT���� A��� >�����X�{t�F8\�l� �?��Ңg0��Q*��v��X����2���]���D�}����,?�|��<�b����I�O��ٮ�)!!��]x�(2���ү�.�ћq�˦h!M�ö�ٝ��sc0�W3Cx(�瓚'���&;�a/����[66@�%S�_�I�ы3I�̫#b�_2�>\]l������%g��4��*��*7~�����*�� ~��9t��ϧ���!⦒�CE�s�V�vUy�I�3��<L�4�ߥ��8��D����u)Sݬ�}_;R^dH��S������Gb��@)ܹfk�{��G?rƄ?��$�V�# ���wq�9[%L����tz���~��z�dò��Iq�i#5?\����~V����Q�]Z�/��9�J�s?3�-'!!6B�qē/��P������o'r@��Kތ���� �KX��N.���EBО���K�!�KǏ���+0� ����D�h����~�,{4�9h؄���ٳH<���ۋ0#F}pP�#�]w�D����
�ȸ�̌�dSLX0yj����;�-��gk��=;*�HaQd8�#w�����w�Ȭ�9��������Z�'	I��$�r���ր��T?��2"q8��S�ȗl�ܚ��a^��n�S�]��b�)Z�Z�j�-�X�tmx��us$0q�$難��0� O
��X����A��3��f:�CGvJ���/�C
��װ¸)�xs��"��U"ءN�Gx�6x�6�7˯�\���g�/�!�x4t�ߴK%C?7�?z~6A�+�ͪ�AE���\��vk�z�3�;w0k�ɣOa�=O�⒤H�d���-���[BV���t{Ԣ+�b�F������]:��ծ+���ߡf/�i,2��5�}�H������ޮj�m��i�6'�I���o| �FtCs�_
N3y �~���As�uRz��L6�#�IT�~�5�R�ߤ�! iM��2Ǔ�=�`B8�
ȃ;��r��r��6tK��Q`�;��_�}J)��3�Bpm<�=EQ��|\$��K;�$�kvfa�{E-�)j�y�O,��,~�8K!��|#��U�}*[�ͽɎ+y�!��<��=��^��\�����a�dY ����ؿ2�n�w��4=(Z���U{۪��Lb!��3���V��_�`D�aJ�!b�Q�U����[��8�)��e	�X/�οl;�T}�-U�6<U���D����J�B���<�JW؍A�ޑ�o�nf���W���_��MĤ�Y^��ϗC�T�Gք�Z{W�yv�I6D��6�$���[`b�� ���Q���G�j�4A1.������?�q��C����}�L�(���4�Z8�/Y��e�$t����xc��6�L��e|	yN\�8qn^�^�;!m�L}�w^|��(DˀAYPȾ<~��ii�wu>�˭��:��6{��ɣ�����>��c���e�㐬M����tfUYsR�#v����N�W��[Ƥ���M�6a�c���ԋlo�[m�G!�	v� T��ZE�#٤W(  �v��I�x�>$`_�s��J��:�@%�O�b`K��v()K��i+�?A��<��bw5�E��ճ���_֣��״٢�[�/O�l���8<�}(�Y�H�mO	f=4���DA��cb�2$��?1���d>7֊�b�J��O.A+�{�gJ�/�4<ځ�g,1�hN��m��c�/R�c�L���1�B�N��rn��62�n�k�̶nk���L�.���ԥ/T��5b���}i�=��a;�������le��U*�iտ*�B~��\�6���J^�!WjB���]>�t���/ŧ�G��6L�T:c�7����5_��=.Y���c�՟��_�>s���WR8:[o����J�^� ]�7d0:���oE^����!�;m��*���л.ַ+��E�m��K��p��S�N��SYܴ��G��^7'si�3���g.r"��q>.��\�f��,���Ʈ񥯟�{����pz!����G0'Ok/��/I���pu	'5����+Ϟ�Ĝ���"��c'�1�B��7htr�2"6��v���r"7h���|����@YJ6Qm/�#������h��@c���;��OkE`}i�ז�8-Ȝ��!:�p�^G��(�b?����E]->����Ű؏��B��%�L<�/�����d�*�-�QC�4PT&�Yɱ�u(x��~� 8@)S��vD��^h���Po�����W� �>T�	��4���n��V�R���Խ�Rd�n��Y e!��Q,s�Z�%��i�>R,{�H$!�z�@�AhZ�<{��k�=�y�S��$�d":��=o�j$Nc��^�mg�u �hj�s؉�r���Ԯݛ.y�� ^�y9d x���߹�e��˴�oo�����\~�[�i�ƚ�'��s~�\KAe8^�ɪxL)8�Ǥ��$�7��=�<z��8y2/�q��]�C���(��T�0W�C&t�-p����{p�(���TP%\�eW-� ���j���K��ȒQ*���&j<=�0�m]���_� ��_I^u�Qw:�|$�И�֧:���	�㷽�/�m�z�q;Qz�Y�ӟu��>j&[��/ņA!��؏�_�ڕպY�X����c{;W�-�S�k���Lx�F��h�r Ï%3�6��M�:����4�hO�{��ֳ���#�Nϋ��<E���Z�M�fa��W��}�J��~�����n`��pU�2�/�����iF��*֗֓;�;�J8�}x'΢Ykxx �rI�)��`�_ye� ǆX_�YE���l�B��5��%oڅ;�k��öCv�4_P�L�.sAy�k�7�0{��Bڮa���g� �Cĳ����\�͛G�N���@��Q�nhjSc���i�5����Co�J�4��N�����=��"Z�����D��<�t]��[:���á���������
�u��H�5z���Tg!���-3yj@�:Z������>n�����̑��`U����IdJ�����1����8#.�E�`c��j:a�Ƣ���7��5x��@)\)K��]9�(��>��x��z�LQ���㗸�l8�֗��	�J���}츯"	h��`%}�6����N2��G!+�SH#[j�ϲ��:Z����ڸ$,HB�63�~�(����
�f7�A��L��Nޕ�:���C��erz2ۤ�����6�&�"_�l�e4�k��jϯNq+S��օ��"�'�f��~�qֱ�����\�x^� ��`'�N����~�k	M�!�p$$�qh���g��GtH�`^w%���3i���{Z�$��'��7����9�{�����:	�m&��CkqX�)�H@Fh��u��7�G�K�pP�]h��tP�v�j��K�2�6��3�D�}��Q������o$f���#�x@;d��v�m�XC�A���ಡLc۝N�'L��Un��S�#k���1R����M5�nE�k���h�q�Ƨ�K�<R�o�m���M�d$�K�;1����U,!�|'��n��F�
wg*˦\����X�N(?�z�MJ�FA�����t�ڄGБ/���h��I��.N%�D�:ƾ�T��rcJ1��69��J�LK���+�8�}|[z4aJ�����������ޕA�#
խ�G:�欙x��3�{{Kq}b�Ij�|`��n�@Zg����@�}�^,c菫�e�dY!����o��E*t���\��A �<Cuo�'�@5ɍ>���340�j�9�B[��tT�-l�+�V6���9P/fD:�)}��|��/�\^�/]��-�æ���NfF�|~&�Ո&���+5d�m��������NL����7�q?����� �K�,r�=����u
��K�A��`�]u������]�a	���xs�	Q;���v�q"�B.b{'gU/c; T׾	�	�h�����F�-
�D���@��_,�;q�B�[�w���<­��������ri�<�̈́
;�ڿ��aI� ��-�浵�xs=j`�-��&���R
��Ii���M��+'Y׏���+�$�~=t%��]�`,;[��ˍx�c��)�\�3Ӳ)����K�b>}��̚�l�{�f��,�c��a�L�}}<2:t�J� �����f�t��9L�Qf��ʭq~�P�rr ��-����hr��nr�rD(|j�Y��V���Oh5�Մ$�Ba�x�
6�j>�T�����R���K�^���O�!���ۜ��Kugs�����#r�m�r)����Z���!|?������\u��=�������c�\�%��>5"N��`��fB������b%|�K6eNj%��`�*�mNo4�`�]ƒ����Ux�v�1����\��W{_�[�m���'���5tʢm�"���灅���@R� Vn�?���OJ�%b���*�������l �h�Q}Ӯ�E��6�R>Y������b�gY������hy�C�!щ�/k�/�3$�1��=�QEd	�h�VȾA�Q����͒����'
"{ύe��ӫ^[����Ǭ]TJ�B�zQ.����Xe�.��un��w��:�QB?^@�Ch�ȍ��H���Xtd�*�>�2��(Ma��x��Sqxo���2����6���1��aI�o3lW�s9��av��o�R=��w��$QT3��(}/�q'<�2�2���D��J1�!�R�x�R���ZA��c�J	rHC�Q~ְT�O}�bRorx#���,�	� �;�K�9�v�����D��*���7L��=~������DiM��T{K���R�����A >��7�cehׁ��7�C�y�p��}!�%��w��8;����]�����C����1���D�h�j�Jr���l�&�C����)#�׈�r�a~��2����i�������K��ٲ66�\d�7�Fy^fXd��&�y�W��4Tɢ�<��w��>\Zxߓ�͵_�{���X&��xm����1��X��Ia�8�D�/�* y��'�gg�Z�UJ�zm4�Z����H�N4($�����-J�b�O��������,3�k�$B�Ύ%x3�
.��R����٫*�~�+5�
d���%tƂa�������)Ӝ��z�YZԈn��^>�R�KD��nl���؞Ѱ*Uv�wx�����_�^zh�~��?�����l6Ñk_���C�:���bק[�+���L��Fv���F/��80�n��di���5o'F��߷ 9�A�J��~_�\(D����[Z�t*��e֍�^����ʉ+1<�Q�5c���@�� �~���h ������z�}dZ �!�.��C[��(����N��"1��P��$�!���0�hdKL擄P൏8-���L}��S�琏�e�[�_��G���CH�t:�zjL��Y8/W���p�'u�t`J9ͤK�()��ZU��q@>�R�Y��~-_6�fO�FR�7��m�-��D[��#�:�0f�l�`�(r8[z��U�
~�.��֕����Gя��V��3��B�S1��{���1�V:���U�po�)��Ċ�%�2�:��ЎJ�j���̣M�i�i�\7��ctȻ���������?�gϏ$�և�Qb��ݔz\�7�yTg�6�,B�=n��S��B�>^N.�_�����
p�{U$s�}�pֹ:8��ӕ��X�����V��dlsm����a�#����I&�Y����a+s�ò�Cne2����{�gm$���|x�ϲX���N$�6���?�?�^�%Fn�:��aE���Y_Լ����F�e4���Ad���������,*���s�%���{�M��I�t���$H�}�
��˯]�{$h]r3�n�{q�g\�l\x\;�^NQp��е����g�#9E�MT���,ɶ�U����V#��~7�z��?&Џ��Y?�c�r�=�m{fZ����W�UͿC��{sp�s�:��N)�wP��s�A�<ͧ	qi��ZM�
Bج�Gk�fok��Ӡ��On�/�8H/{�,|,2l����۳0�b�O��C�G�'ۇ1�s��8�k�[�wQ�9�s�CVV���;��7�8���W3�[��׶e�2����:.Ґd�_���E����B�s6�RD�>�fB������I����m���&�ލ���i���q͛�� ���Փ������ ���U;��ڲ�����R�/�l��[����F`�ʳ���_����JV����X��=���z��d(J0�$���.E^Y�Z2UR��=������x����q"���\��"���Ǻ�P��1��zAWSE��\��=<�=W����7�M�jBqD�E��<�-�2�(2�p��\��5"X�J�~aV���O��/F�����Y���6_~?�ԃ���a��ZDy)!SO�ק%�Bp����w�X�92͎��ka��a5�?o�2�R'�hh��ۙ��[2�H��1�?���M�%Oc;x�t�]�U4c񶰼]��O�w����M��]�<�z�t㠬�w���h��E�|գr'c}>��EGƄ���-+���/�AdgöEZUd`�Ƹ�
��UR)����5Ul-�|�<�����*����{]���%֥R��
	�T�=���#��p��˺��07e{�K��Mj����]�P=��M�{�_��r&78�PyV��� ]L�uIɓL���u�kǔ����y���a��������C�Ez���ۗ���!�F�o����,�Gw���IE1 &�������N�B��3B����(�Q[w�S��u���b�?ɣ�s=3���b�
��hY!�CA&��j���m�	��dV��&f�Ii�ᚼ$'\������=�a�������'<�O�p�Քћ�Q�����aP:�)T*-|'^j��n��D.2���v�K���r��Y�*Vِc�<5����JҊ�2�h�hr5��3��0l����Sq���l����[pU��㒟_�q�t���)����=w�tnR��m�0��菽":�FI����a�Q� �w��h���3ϳOb��@3yԟ������fqL洽���Ľ���뒪��Q.l��^x�0\�ٔKsy�[���b��D&����e�����hV�k��L�2�BNm��bΡ�O�u���g�4`�X�O��E��"�͂�׮���fd�U��g�lI�}�Ch��HMH��anc��[QQ���|�h�+Ԍ�RG7�ҳ���#���EpC�T7J#�p���4��+9l�es�j���K�e�Z-V&7�lGہG]e1��~���;�e�ϚXA��\�Z���.�"74����`k����i���XNW%�cg���a-��I�K��R��w�e����+�����5�O$��z��!:����#���)efQ����S�#������Ż�ࠦ�Q�EW������H�2�mf�����7i�K�)��y���&��iY�	k��~�v#2^�G+���2������{ݍ��@rQ�����B���&hu������j*��ΐ̀��2� V�O��MBT�b�����^n+��7:TT�*>�n�t�֜�y��cG(���$�[fn��i���.�o���eO��6��͌T0��r��7�Њ�7Y	�ب5yh[�Afm�#���x�f%��
���k8F2ך�1͍�rV?�Y��4��u��M-p$�`+���Z�x�(�*&���ޯ�n��<*���x��A���]�b;+n���nX��K��K�L�l�t�,����k�x�j���>�׶��z�2�l,~$�Y-K"86J� �ue	8�~�n����B�b�- ��J�����N�[�gI@햿�"r�2s�E�8F�7���1�/��\e�� 5�D�&O��0��=ˢ�N���T]�&�j&��Cv&�O�8-E�T�s�
��x9�r}N�&)�H�����K��I���<�+��5O�����{��,�a��k���yq��,q��1��w����B&?�Ҭ����/f�jzT��d���=-k}�Q
�O��B��uA���&c�<�}��c�s�"�%C�K������#e-���|zvL+��\n��mNm�݆��Uda��-�x곅��Τ��)f��"��5v��2���U��Q�SL��I�'=�RD��%�d��{��4Ok��uk��K�e��xĆ�������QuՋ��5�w+\:�J��GeJ���.��,l�~�A�'m���*��)��+"T
���%ѻ'��ĄͶ��֘x���g���!�H�ß��4B'<��tu�K����'�Ѿ��Ѷ��L�1��m�9Մ����2�	��l��w'J@�u�O�~�	�[H�*��VF�����"�k]S��z�	���u1�X�3�x����
�N��sP�:�ٳg���������d�X뫝Sel��!5ÚWC�8յ�c�Z�,�hlVƋ�J�*�Iz b^�T��6>����b<�z�`6�AOy�O��>�Zp�B��;�����vN�r7�x��*Uh
��s5��F&��d�\���n{-��Aڋ<��e׎Ǳ3��Ag��$�K_'�Z\���G���$"r�6���>Ӓ+Ǫ��Y��>ɋ�W�*Ü7�@(�)e���Z�@B:��Y"�T~Ϝ4��2�y�|���&�;�.ݶ��KZ:����m�k(�zoaN�[{8]��A{!L���˂>���hq=��K����sk'*���!�O�:��6_\l͜ac�r"��S]�8��ظ�ӭL�\8���g�>�șd�a�N�!��=�a��C���n��f�$����kv�_n��dc�s�w#C��}�a{�{�h���n<�?S�xP#6�	�i��q9ݥ�Q��h��6%΁w�U��,
�Gg��U�j�l��	4�=�E�z𑎾�z�8�Cu,�;>�����v�)X�hr�Cر׽|c����?�C]S��ȱ����y����
{�zY�$	��W �Z��-��>�k�����ֶ���>�ڶ��a.U���Grwo)��
Ώ��(9�����Ǜd{�����/��[z��4g��,jk�@\��L͏y���#Gd��
�5l9���Z�^�J`��0	M"��L��H�Q�$z��/�+��z�.v̌&(�>cx��f�����7��M؄_�L��1Z@�;���&D(�<t{<i�+؍����b�������ז��Q�F�!�����T|B���z��*����V�*�U�u���G�}��*����	8��w$��~b)W�0�]6��vX����8��Vȅ�{�ED����I\� ���(j�S�p}g�=[���WƇ�
�Z��h$�Y��1Ȉ�x��� !u���-�l5�u8K�>��ÒF��^P8{e�j�*�h8�;ǫ��I5'�{���`�æ�P������2 q�H��Q���,w���@��h����&�HM}2��|1��7eϜ*��蔸� I�^��Ս0��uc��;2��	s�ab���3|�Såù�9=����)��ƕ����8C��C\�輊RI�{[�o���[����o$e�TQ@����+�n�e�$�}w�?��5��K��54<��n��4�wg|RF������')[���c@��B5m�-G*=R� ��۞��)¼��^pY�-W=b�<e���(�^�y�~9��n������k���|tyK/�C˼(���s��t�8��.һ-S��(=�d�z8�攐��Aؠq�s�4�n�\�e�b��h.����R��M"|/ �.U��.�I��4s���/@���6�ZN�#GN��O�3���6�?hc�ͪ]vnF�w'(-3��
�r�Z�u_���J�?f�N�W�.��}?5��ߑG��~�r�S�0�.c(���"3�b�^�t�c�&���0��?t8�\�i2^$��h`���T�{q�Rn�$ťg�3�؇I���ve[�./�������23AS��R�iُ����K���AW?Т�ۻ� �r��m� �u�/w�B���D�+�Q����!��Z��Y;E��9��S�)��)�BJŭ��dPR�g`U��h�ٯG����o��Q;Cn��ZU4^�Ȁ6�AN�]b�Q�.sp(�"��ԓI2u�DMM�����a���c�|��P?P����l c�x) ��.���n��ڴ8y���b@5	�! �D4|����<�ɰ�����h���<�� g��'���)2���S����Z N� ���K�k�D[�n��`�G�٬��v�Wh�Dk���:9��e/�ן��B�Z ��P3̵�I�d>곢�3	)������|��"�m�y�� �k�Od� �g
�X��j!��V�GE%ܧL��J`���[�w�{��׍#���K����7:,("�2z��k8O%l��j򌾨����E)��{�/��!s�x{�(.fz�QH��oF�K�u�m�2ӑ9 �����w�|�nQ!�A
��7�ݩi��T�:,�fOqVς��z;f`Jq����
�Yw.���ȸ����[(��4�w��M�=�q���Wr��g��+�ju@1R��ʦ�u=`b<�˓r�B'��~e4�e8:�rd��w��d�儹8��At9�S�	#�W6��L:ec I�覩κ��Ѫ�o�]
�6h�ؾ����� xNmV��� �{��~�*��^r.��<$�*j��谼;1(�5��z�q4g	p~iP���cq����c��W``�[�k�����d��{	qp|�XȜP�iz��e�]�-C�_P�Oϳre��ʹ�Ml���0�����*��N��UѼa��;(Γ���Jo^��������҂_�Hg	UAQ3�m���_���>
���s�a�#����'�/8ᗘ�7:���e�^��%voK�Ta�[�M)'ȧ���봱�����8S\�W4��934��n�"�ۊɲ6+ղ/���/+{pa��8�	YD��z]U��
�0������~K���<����!i��|������,q�����B�d��W5�$rmNY_TAvCt�X�5��mK���>��`��>��`�����El�����d$W����D'����T����0G�"�6^\4�c�b�g�,Y}׽��CXj{<�&=k�Y�Ƶ��ѻ��8̆�_�7Q��P�<�c_�c��#����j�e	���b�y Xo+�E���T
~wp�������'�әn��m��>��-fl��/I��ݚ�R�v��]&9��K�b|[�"V�O�|O��D]ܓ|�٣�yP/�� [�Z��iǾ�a��Q�R�$��f�[R�l��}_YT�Ph;��:ܹ(z��g%���q�e�������������r/UnTn�Zs���~�3�d93�E֧L6:j�l�E���%�(6���Q�Ҋ����f�k��� �����>�:d��XKt,��f,��*�*�D.�؎�0�
�88�^Yԓ��r)}XƓ9&[,tV �˻�6�<�{��󒝎@I7j�]���f"G�w)bӲ�Az�ִ��є��������.��`��>�6�>[�=�j��|"�I��	��!W��}Ӷ,%��>`�����'�#�#�U�Ƕsw�ؕ}�$�r���2$����Ų�O>���]
�'өQ��/ҿo����#;���Ѭ��������P�����[� ?.��������~�Z��\BA,�*rq������ڬ?z}"�S��m8����u_���(*����4H]"��%H��!�RR���C�#  ݠ4CI��~G�Z��p�}��<p�o�������y����-��ѾHd�x�U(A��'/P��i?9�ȇ᭾I���mQp��랉ݏI"�d�z%��zi������혫�y�N����H�r@�:�
r��6��;�Z��bL2��;~}2�Yy�\Q����k��-��J�Xd����c����D��6�t�����$6�GR��/�f��b#<���և-��V�&�jsInn�~�E�L�=�� -E�72�H�ُ��T��\�L���e9�u��o�[I��I����4~4�Of�4R��k59z�@P�����|���Z���wI�*���u)��"��!�!#^��Xj75�J]wp��CԂp=u�/6�f��_Ҽ�<m�:~��η2c�Z-�حh��ަ�JB��=2Y���-��>p�T�ſ��E���K�	4n�Lq9:���P*E�;3�x���X,�r>f?;RPћ��N֟�n w��u�|D{p�c�z̉���d+�\�B���竆)ep&���Y(�N��dz
#��9���ϖrG0�T�CW��ص|��J�{�:yc,l��d]�ģk;��$oh�J�5^�W=ɳ�	jH�o4��x8�\����&��.���$�2dsƳ�Pٿg���۩P��v��rš�W�9?�Z���7yZ��!����9���*�m������	���/�l�_L"L�Q#F#:����Q�L}�Ɲr�|/�D�a�ј���Б���m���H"T�;l�ёϩ\ι����O�*R�j���H�:ˡs�X&EoB>��ٜ�nX�xS�د�!����⸟��������vq�e�� Ș�gq���"p$�ˮ�`u�K���cg��d�� ��i���<J����:|9�׬1����@k)^��U�%�#�G�F� �	�j��Ϟ��	��u�G�s<�״�h�����k�9G7�?�'�v����\Ƒ}p�E��ф��,��|��s��)��=*�kY?�b�y�x���W94�|��9^��y�S�u��q��Qg�CAA�f�C�Vo"?h (�x5�\y��,\�x��XP�� k?{Z���K�)�U��WG���>��c���]!+���No甧(z��ϣ���بh4��0,TQ�x�(}wyhiuÞze��u�Ӛ�k[�2�9F�^��'��vq�/�Tֳ>�U@�z�5n�m\�E�2<T�t�z����$[���������l)J(�	> 3��pu8vj,hx��&�_�Y�F�/ɳx~{�Z�2���>��1n��)T�~�Z���"n��@,}�'�(��^޻=c��x.��W3�_p2�+E���CL8Q�~]i�O/�-5NEG�>##J�J�#�$V��	B:�*f��P26�SU禣7�G�,�����!�c	����N�;�+�š������2����ǭ�5qTW"�s�K'��&O�q��ۖg�dVC���L��LL���O-���53��b���i�����BV��^���~��OH��P�^���qz�� ��	����i�@7M>|���)H�*F	��ry]#&rh�.ڤ����k���u����{��^Ц�@�m����)��!�j��jY�.(zkB��u�}!�=��R���q�*A_z�}g"4
)$�C ��h�Y7)�����
ə$��y5�zE��Е�L���r�"�V���:Q�ݕ�����U(=}��zc��׎0��sg<keS�!��NfRo�M�mbY;k��e���5�z�s��q�E�������u07���7���~����1��ώ�_�%���25M�2�Ɨ�����$�U6g*eU]�p�#�IX�&�%I��tZ���{����[�k�'OVJ����筕�'���ߙ��$/�������te�,K�B�S���*�����S�����p�?34N��q.�e{h�FB�>Sr�i�U��mu��mzK��2M0ځ�v��8�\9��ㅖ?5�4 ��h�/8ҵb�a#╌g����_a�U��Q��WSѧ�6���J��'l7�`"��J�0VM�,d����:0� `h�!:px����/ZC��?1�PS�BR�ƌ2�@�5pr����|g��Tx]gQ��Q]~���r@�q�dc�̛o$�H�ӟ��O�κ8&mx���H�f��Lv�8N��:��䶋�A}����q�ۻ�:ڡ\�H^����eH��<�x����>�z%M;���*���5&1ڜ�5R��űa�5sb~��|�[o��iP�������%q��9o�gG-��JЀ�ko@���5�@��s�r�!rcVJ����õ�D�d_�A�!���z��˻;j@�_<`�ܐc��i��@�3�Y4��c�	<�ʂ\l�*3U�ִ��;!@�|)<�z\��Xb��L��%������1�����]|r�������l��le̟HmŢP{X0��Q6�%� ��ǜ!�L��4����q��~7�(��Q5�ei��<����=�^^�����&5�2�G��[�B3Q�Lc������CH���3����{�h��×��s�J��L·�c=����B�"�H?zN��M:)���l�|r�o<��f�C�S���f<WL��ģ�G0`mj=2gHI�F��u��#��;��!~y��&�?�Ď��� >��$�IC�V�X����S3Ü4dў�,��w3@�b$"��e�ó�cakY�kdȮTm��´�������>�iя�*m���I��{c�:s��:^]�-y��������*�DA��v��!�v*�k��&Y��J�>r�c"�<��3#k�/��Z�S�^��pM�kN<�Yjȓ��G[���M�4��>-Z�[gn,Af�L�dx�cԀ��l.JB������}^#�)o��Y�g�1%�.�xY�o^J�a�ޘӇMĵLG�+�];�I�+���y����u���u���`xw��I�v��P_��^w�3��&z��Lϓ�x]]�n��o��'Az����ʌ65.+�6CG���s-��}��x���ۦ�.�kf1Jj;���圌s��_���i�ڙ����t����u/�k�Y��S��q�/ܷ��٬Z��т~��íM���&�-�|� ��;bI���x�m���K�P�Q�ʝ$��l��-�@K���;<(&�5TX���ɞ5�~�?��x�?���q�P��8���_�e#XԶ>\�\8�/x-��9��hB߭���p[@����R���h4 ��INM�q�i6�&�bZ���+�'���� �J8���Ir*�Pu4ө�`�5i�Z�� �S<j"�r��}�ņ&�f�Y�������!��%�	
�+շg"�>w�
�.���+�Z�񺏣y0G��#/�(N�q�8�E�"+2��Oc�8k����ΐ2x�kW׉s��I!�}�ͨ	�^
m;�����u=���jFǅ��/z��a���%H+�E="�6y-N���'�� !`<����$��4���~��{r�/����ce+��J�&'��z�K}>��X�6?�a��}�=Mϲ��cz-���$o� #��d�-P���'�V�|f�~���誒���ҿkd�G}8����>څj��&u]?Z�Q����3�(�_��6^���d�E��gz7Sg�L�5���������Z
�����&���Z�}�^���T�a�a��n۵��Y�z��T]�֏(9��������)��V�z{v�w�ڞ�6	�?��R�]�u59y�T��Ae������zƂ�B�Y��p��P��sW�Q����A�����Ec�)E�D����y����$�9�����]���յ��t���}�O 3���G��F�2AW�2ym�yG���?׶�0y\-V���՞ ��ɳ8XR�e��:r1�č;�*��&��v<�&��V6�X���k�%4t�`�k׷����ͪ�[��QAf�_�sf�"�԰���t��Å�6_�d���B�V���W%�D���F� -4��
���=b��k|U=��v'�~v�DAq���UǾf����`�����R/e�=��'������W+Q�{����Ѳ��^��	q͙5�f��e��l�;����u�-m�b�|nj=�bc� &y����r�:Q:�W�/A�j�NZ��w�!]u\�D�\��"/!��}�Ŀ����ޠ�ݴS��:���#����&Z��~��<{�x\pe��#�I�c�RF�a �y�H�J���V�B0�PF(;Yc]�~����˃��<0�lO�Ŭse�NO�n<j�Td�M��W��;�s~8f��9��9^M ���N�WT�tL� ����y3�)$l3����G$8�}ڄ��!v��3H�W����>}'�%����eH��+_�g Y�T��H�������AS��j$�|ܱ��w�ԇ��Q;�lP�1铌�^����͖z}w@$�7�(z�
�M�U_���(���
z6({�5h;��1�M��c�Sz�Z3�;�"��[<�GF��k��O9�FZȉ��.��c_��n�5%h旋��0� �0�r&��(����-�k�Yd�7�8vZ�h#>�1^�,
s`�rit37�;���u�M�8t��X���F¹;9u�;9w���9��������'�]�ӧDx���w[�"P�c7��Y'7�\ܝa��{�����틓�k`�j?�S�ר{�PA2�Vzn�X���A�[8�Ԗ3st���Uwl��4��˦r�w��0n[c�޳�|t#�~j�;3��9�Y9�VJ���=Ӱ�����"&���V|]NW�b~�L0f(�>l�Vn��}�'��%3OIIkor�㼓�Fy��B|q"��}����D�i$u����٪'��z��a(�
�&2�čT����<ygKDk3�M�j��rY�#��F�^����tc�n+:�&�:-�����G�զح+��؅�X�x<t��%]�%XY(j��/�&3o}o�5�LS��&��<����_�F\{;���v3Z"�܉O��8��!0��݂�Mh<��;�p{wD�9�9���P�i'S]pÏ��	�&����\%�Z�x�
��� z����yS)z�gj0��B����f&�Ou+D�ƳV{H�rB���wd��Pj�G�|}P�ݗ�/c��ӆ�8@x�3	��#��y���r�����|W��S��U?5
�}4�.�Ϡ�b����D|�1\�b������"t���c�K�de"_gV?�QSM�W���qV;�Uof����~}c7bT��w8�����I�D"p�|N<&kW����ɾ���	��_���t���(M|M��|�@gG�9��;=��8��W�x�uy�� yUZ�'WS�Gu-�\^��[�ߣ!��_'��bz�se��h^���1Ĕ�108�6W#�<��9N=C�� .t9����+����O��Y�d�#ܺ��n~Yߢ�I�r�����,��J�IG��N���E�{�d3�̄p���}�+�c����i��Тk9ȸ���c�B����VٜM 7+���t��Of�ii����*��~rp�Bz;#�]u�<�*J��}���!���H�]6��q��],��?����0��˱����QUT��$��}�"��C˻'�<\��8{�?��LdPSW-��	t	���y7u���p�r�{�9��	8����H��,9��c����$<<�ErK*duh#�(څȔ��9����U����x��_���Q �/(z�xL��H�O�WHz��7��dv�e�rl�����Emլ�	ʒ�Y4<U2h`�O:���(�D��ZЈ��ϑg7Չ?iظ&��L.Y�e;��M 6]����s6��AQV���Z��{L^ R�jr�{�N h�n�:�����e�;;�ą8w��'y4���Hi���ź��|�>{��;��}5���U�ة�V\��H�#Ԫ� Jn�uYV��*>�E��dر��*�~�~[[GX���sՇ�J�W?H��{���R&���e�R����uS���?^��p��(���I@�{�wJ2"�Z:6CК��|5�)�W�7��/f}���H
?AV��	\^ql�.���v���8�9	?�����ǳ
�����;�����ٛ��GP&�7�I�/�{!��MDA|���OZ�A@U~uW^���.����q��࠶���]J��pwQzVa�g�cTu�zC��*:�%�����$�:�����>�rshI6��]���5�Fv�Z�'��,�h^F9����ps.j�>�MT��شБ�`�v��!���6�zJ���r'�r��Ȧ��w�z7�d��`���r̫�Ӥ&M��V��q�'"��v.�TH�b��K��kx��.����Ţ���!��� �Y��GR[��]��-Ԍ�F�Ǩ�E��`��{��r=���f��]hue~yK��|HI1��=g�.�Z�?*j�G�6y�*��<c�*��0����p�:y#|���V�yZ6%E�U&�e��[��/dje�8����>?��o�?�8٧�5YDRq�?�R%�aE�+0�de؛Fb���E�og�L0i���P�ǺXX�Vz�J�;�Li��2�Ů�/p��tOR�O3�G������h��Ox��6��*�E�r�F)�ո�[�GS�$�H"���s��(��<f��"��Y���F���o�#�2�t]�9�q�!��+��ˆ���D/~~T�"�c�Tiڮ�n�PB��T+	(�37�Ƕ�D��ża��q�I}���M�����B���1Q���C������;Q4Y��C����ے^�Y��Ӈju��>�Dc�f�w��8�Yꃌ������q�X!S�Ķ[�A���A������v�Ł8�U`��<c���uf__߼��~��aBwv{;
Il�H+��i8�^6�d5��c��B9�䰉CV?��o;����j) (�VVa]���̔⦧�F��Py�����}�����Ç��b5����~��
��Cm �NR��Qݫ ���[�vdX���)�K5�H�h��!�ԩZ$Q
���φT��>��r�L�e*?�@F��m�x���ȿn}�� ���҉��GX;�]N�m�,*������ύ����rw�kAp{fd?Y���;gA�p�g��r��j���!��7����� ��b~Yxúb��g�o�X���Y%;����Fp����~�$J��#A6$��QF�P4-��������'�}������LM�����?y�3�FYIʾ���st�P΃$��l$���G+_���#����l ګ�iW�Բy�n�ʢv�x�;}���O�Z�t����l%�b�@������̤��u���?����XV����U�e�ߗ���俼����_�g��a.��j���U�K�>>�23?!�����r$t#Y���D΢�<��L
���|礥�|w�~K�z��	�O�%�uO�O�����a�:�7�\��'ia	��Q�X�u�FU�K�Ců�t�������e@cl�_�H�GL���<I�vqN�rpw*�rvٯ�C#j�o�\ӸS�{�� ���"��~�?3�;�ӭ�j��w�i]�+�^a�ӃRݨ=
���ü�����������c�Z�i���?��tױJ��En9��z{]�����^w�I=��)�?{�O�8o]P�n��1����q�-���+��w�r�?���V�v���|Nz�nv�~�,3ikYpGu�3����3�_��cO�X��!ѳwi����mdc�q�}�a�݂���&�@����[����
I��#X�.���o��T��q�����U�B�|�y��jN�ݛX����O�&B�����J��H��΁iO�8i���vb���Rƪ=��&����u�k=��%�7��������|qh�#���`ކ�?+ֺ�ChWC�g��Z��o���T���w���I�kR����ۈ�̓��3��"�sn��`���0^��g�;��]{�:�9�V?b�����Q]\�^	�Ť��;�]b[GnS�#�:$2���"�O)n���Z�,gQQQ~.MLa�PL���������n�`�S�4
�*��K-f�����av~e%��W�Q����O��:]��SR>�0�����J�����?]�ru�1}��5c5~�r���>j焐�46WH�&�_(�����oaoz�^�Л~�+�ù._V�64�Zm�5ܴyl&��-��s]��J��u'u'�{�����h��R�|��MJTxx����,e�3Y�xѡd�"��Zz{&-��_2{��ϼs�����k~�3����;z�iZ�
�Xff&����X���Ϥ��Bȳ�+9��?,x9��>������L�(\��9y�9͙�GS�v�$�w&�TX��Al�v�X���^%[���r�cdd�\�zL��w�Ҁ1[g��!Z�aLSG��E�}+H���X���w#'�3d���~ێ���D����?;�}+(j֎��xC�irI��e/���N���l,�1���f�Ճ����~ҹNȮm����
�~6���#�n�ۄ�An����%B��v2���Й���/�KG(y�>6�a�ų��A��:��}u��!�i�;(���7���E��-˙����^�m��R��zWo��Z�)ZE���_~��?�38�	̥9zzuu����ݨBuEی�hc`ч���k�,`o݃5�wǷ��^���_�3�IU�gZWO_��IW���ҽ���%�J����ڒ:ъwL�ο6��%�A�ya��e��wd~>쫲�oNң]t��1�x�\c��ӌ�c��k�Mz^���ϒ8�=��q�Y����DSN=��)�fj#�]T��s��h� $���E�R�I������ۂ&FFF壮�H%eeYq��������ȱ(M�w�}���#�߂���2�L۷�y��Y|�W-���睸Ӡ��gNk�-ߋ��m�t�Pݣ�db�� ˿�#\� %k2o�Ĕ>�".�Zp���ƚ��{hs��t|$�Ժ�Thj����.�x�;�5]��c��x&ߟ��p���4�o�"����C&w��
����%�����-\�=�Aڝ��k�b�b|!^�F���N��>��Y&(�����@�*e4ס������닏õ�jU����N{K���<�H���ӆ�מ�K�/��>V�.;��oe9�5���#��;݇��&J��Q��Oc�
Jf��������\�ꯢW�k��?�N�'TAq{.~�v��@+&)����pz~�٭Aq�O)P�z�xF�i$Ƕ���HuF����&�^�]�͙�FȮ�P�����*C��M@��Wh�����XS�\�Զ����՛Ivp<�E_�피�f2s����dvH�������W��2z����|P�v�h��3@�{[�lI���t6�E�u�z�B��4�%���s<{�Xk����������c�����{���y��\�>��[q���d�4�{y����-w�q��jm�LL���5�E����V���y�4?�:���Y*�Ly�¤�mÃ��$^x:���%�ވ"i5�i�oq ��{��x��#�
����a��f����ҹ	g���#C�E���f�z��N)ـ���|*ާ3n?Y�~���`���U�sZى�/�>x,�oߺ�����W���.�M�g��
��S��'y���_*��M�ǹ=�}zcR.�s��J�j�@�!����UM�9��3��L,��ް-3k����(��PBn;p�t�9�FΜ�Y�\x��]ݙ����?S��V�k��qwQ���S�7�᫂��{�ˌ{�$��o4xO,� �$V�:�R�eW����f��j�������_���ay�������Q1�䰺X�ұ�m���3cb�qi�t��f��vH �̅bי�LS���7�P.��KA��'��z��Xx��%�7xiL�����'"W���������*�X��=�:��˩,GE49�ɨ��N�G،�Vv���L�[�K�0�I�ƵU����Q�h��>Y�æq��K{�A?�4�+=L�Oc�3M����g!;�ܒ�+�c��5�3��wZ�`�8��ƈk9(wǻ"j�՞��qe�G/�.�<>��lrݩ�{���.���\U�ś�3���[��<ns����ٚ�4�M�2N�_�r�o�.����p1�Esm����(;�]��b!������-4�1�y<go�Dzy>X�ZoR�wϓ�������>y{�;ɬz�tv�O��_K��=B��Mo��X�{5{ޣ�ϩӅ�]{���K}լs����-+z�Ne�$lnJ��8F���|x���o_�]F�N��O6��y��!����N���x�=H��=�~��.��/����q�;���\$[u���Iv�K��n����F{:�*��o�B�!�����3�H�Qc�3_O`/Ϥ�ƕZe��B��&��{y5TG�C�o�]��7���g�㒣������o�R`:�Z�7ʵ��Ef�dί8��u�"�K˴����X.`�Os��@v�0$�l�p�P�d:z��)����X�S����P��ťc�˲�����]Z8����m��Y�^����xo96����y����NW2�,DәfN8Dfk7�E����v�ԇ,�O�mR�tz�̔K[~�����?q�`��8p4rYL��7s�$�z�[�H,lP���@������i#��?�ٶ��]��i[�G���cQ�3.*)K4�5��������Y���Ul4;����
�'Z���G^�Jtnv��t�M&�	��wf����YT6%�Ci|�ß� �{I�g){VG�A�/;߆�K���+s-��=�9��~��])�6<b�w{�c��:\� ����^>��?U���:�J�ѥ�Q�>�V���i¦��^��'c�D��kv>��T�]��	�BdM�a'�a��ޟ���������.nK�0�����2�Ư_�,�L����j�ٓ�w`�|�Q�z0�=��R�ZYLj3ՠvZ�^./9m*�>C�Oi2{�s���.^�7��L5°y=U�~�597�dڣ��#�l��x��ʆ���xu��4KW8������4�>�f�N `���R��S�0�{�b7rhmp�H��*_MQ�ؽW�t�e��ׂK��.�����Yջ(r��gR���rGL�E�}3_>h1���@�i-/>l����/��V^|��E�&�'|2�òҧ�O���
�l�������WdW
-E����`_R�?$8�k����໕;��͚ũ3W�hj'>d���>�܁�j�f;�D;4�3M�9�u��^hy�{&�X\��9��^�Mmn�����\=s+�_�f>в�Qv�'�A�;C��8ά@c߬-��"$��C�4�����������Y٠��k	���I,����6��5}�?V�6���?皝Si�;�p�X�	虑��V��W�;gEu�Z0��E�wv���.,T�0C�a�i�������E�7�x+l�f�K}�q�Jt��$��OTk#":�l<��G��i�xp<)��$��.d}"�v&uuA���u*m�>
��3�i�ٌ4,�{�w�=�q�ӺO���Ю�6�N��N|N+>�n���\HC�;b���c�˼{������µʎ9t<X��.R%���Cpl�7�	g?�tP F�e(����F�����U�mcg�0���U��pQ��9!�� �_Ы0�N�X絩�"e�|��2�~9����tƈ�(���<E�@ĞxUL�1���m}w�[*�x�$�Cbk9:�*�̕	��>����>�z����Y��Pdl�sW^���[��P� k��%}w�i��e���E�Ӝ�PKC:�?��0�fY��D$}�`4�I4i���	�����0LC�h�S��<~gO+t��N�ՙeJCg����3��Mɛ���e�.�<��7�%��F:��.%:n[�v�uJ=���|�܂�>?�Ы���:Ie`�h��&<�2������KOЌ�a�$�h=���\�0*�	����Jג��07��y��vإI��G�� $\�r��C�y��&��.^<̧�[�����%S�hn��"+@���I�M��еX��[����GZ���H����~��|���螀��i׺����g�H����q�}��0��:�`x��t��?��5�~�V3�^O��֯"�[ ����'/*��m����������=Vu��/�����*�;�&�����Y��;:�5eK��<0O?��2�֣�
�|$�C�0j��.`�f[��x�zO��G��#V-II���v�ᡀX��2D���!�<I����_�f]y��<�"��b�Oa��q?X�A.>����'� }*�������s�h?Y�2h纄7%����75O�����D/rba7��Ε��*�ԋ�*�i:�t��Y�q�N���w��h{z6�i��Y+ڈ��m���W�p/����!87훍}�G�x�$���r���A��j��_%X�.=D/�MGq@���XJ�}�W���jV�4�ĝ�W!�]�7JH'�S&�0E�����q8 Ȯ��aȢ�l[`&����� ˬ^W|4\ۂGL���$�y�,�8؍��D�)���L�+4�Q�ܙ�F&��{/m�rD-k��u�J�W�t�U;���h���h#��p��i�f�汯�,��
�G�?�ɁH;���?A��
�@?y�]o��2l����wC7���V�����b� ��Z��Ul�!%ju�q��Z�Aga�)h��!����PT^n���T8F̷���{�l���6�rw%��o�hh��]��mB؈TT��&�O���#��1���T撩}�l1W������L ���@I��9$ 3��I]83c�������G~xW�F�P�tԆ�Aff��7���[��Mv�
w7���2�-S]PЅ'�=�M��q>Pt@vA0���T�/��~_޺�*�jʒG췧5W'>�Z�O+���QTV,aߌ]�S�8�O�ظ����*r�v�n<K.���Z�2�#]��>1��4����r�C�۷�AJkhj(ǈ���"�/n��斋���۸lx�ö��乵wù% �qW�i�1�B{k�Qk
���1ק��6��P�پ�b��ג�E�������j6��P�,+�@u�K� Kb^��U��_s��j,��nY�a�F
Jco���GE�������'�����t	[u`愈��|��%�%�{ŉ��!��K'�Q{r���7E{�����r Cz�8�����N��dOV�4r�=�}��i���Oɼ���/N{��o�L����<u%`��y��{����+QE��d�{^R��
�c���n��N��t�H4���k���ş%EcJ;B}$�L{��6�L�-�r$�e��<�D�^�R�\z��9�ǿ�7�a�$III��	�s�u$7��=�F���q#�O�/��Qxq����P�p����س�P7s@@ȨވL�s���F��gg�	���D�g1=�ꮣ�ꤰb��Vۉ��>����0�-/o�̃�xݴ���7��4@_Ϸ(V�k/x>vT��ܷ2�NM.h���S�\��_h�פ`��4(T���g����՝��x���<A5�m.�l��A�����r����柟:s�����@�U10k�E��<"�����Զp��Mlç��
�~L��6*� q˒}��Ϥo���m��\dBB�3,�����s@+H����T@y�;�&u��s�66��"A�9q䁡c±t7����}D)�)M*rQK{3�%	��W��ޅm�ܲdC�aeV�7��&<b�4+�_��u�,t^j8�w�	���g$T��c��a�N�zx����ך��������D=�ek�5�������7xypך_4���pU����4;䷮�J}N_�l��u���ᜐ�Gw�����F�sLn�x�:[�a
�z�!�Gy�/��n7��\a�׆�>��;�##ۈASt�\��}�_4G���>�v����9q����gE�Lm�i�0�l#**ލA�ёO��4e3r�����x2	��/�R�����$A��,�U��ެ�����k}z�{�	��ax�$Q�aӿ�PH(���^ֵ˙�����6	��,�"�����INrI�*�� �]6���(Z�J�$�(�э�������cy����4��,1�R���2�Gҩ^;���J�s��x��k�� �_{�X��VRn�Q�i[�߄����ٖ�ܳ.!e�y��A�t���I���H�,9�|�KE��Ծ��&�q����&�S㊬EJ��C���'�xgc�k�\.��j�F��['�=��?/��آh���_����U��}����b�s����R@7ś���
R��/���|�{�ƈD`D�y�����Y`s���\�`"��&q��3L��#��k�yE�āH�*�?z��\+��m����ɭ�B�	������$$4��������nU�@��xm[{o0�Ӎ�UV0�$�ҽ�,+�Hoe�%�	{�NF}e~��RI�a.+�iN����`�}�ˆ�wm�ea*S:�c��^₦7f�#��gUA����z���Ti.L���.�*�K�n�b"�R�Bn�Wy���sj�t�1�)��n"�]��nQ͠
]7){���H���+�N{O��"�!�s���\g��8�5U�U8�P��\&��*wA��"���i	x�-��˼���nt����G����BG`,�d�)�x��Ql��<��������NR�W��G�]��l�^ ��'����xq���Y����gQ�`Ģ4�^Թ���q���>(�wtSZX�*S�h���U�5��%{>�)��|���@N�G�H�Vn�Y1O�z�=s�<�J���a"�<ȨE�(��K��GAAU�^s�@�am0�[ w�ic�@KQ�4��&���iرe� Uf��O|�my+"��ߘo6e��c���+����a�[�E<���-o�T�d�I㌎�@�8X�,��_	1���U�	��
?ӏ��f�׶x�iJ��7MW�9i��x\�nQ^���,Q��P ��x�?�{������$=�Y�7_���Ƒ���5͢|-�y����K.2��b��B�9O��*���1�s敿�ˇ���յ�ep[$E=�I��J=�ʊ���A/L�,l��p�u�c{��=̛���?]��l&J����@nf�O�
�7!��l��U�������>'��)���W5F���$�L������l#��+?{x��P`_i_����o��tR��>�b�7��Y�??��4D���_'���D��N��jz�L�m{����U*[��c(��S���o���:U)�OO4�Z���@+��ݐ'����V��[���W�����$�羃���o�F=��5/l�]�7���ov~��33����[�U�c!�%��NC�U�
�euU�"������7N��4+�9�5۸ZF��hBc��mVz�����a	��:k>�rT��v��A�~�: a��2_sʂ=OP�^8ȧhT����j�>t�4�p�c∺R�2LC>Y�wn+L��I���w��fAs� 5�q���\K_-@PR	$�(�Ag�[���쓖��k�d��&
��rC���\�Icm��׀A��S�����!�P��٥O�����z;~�(9�����@�ʹ����k�1��KÐKGcI�]=�o&�%8z�"����G���΃Y32�9^�������i0T�0)����V9CT��H�4>(1X��#�L���ϳ�{۞�vw7L^~�E�[Z���^�[�}@�_ex�+�vַxG�٥��j�� ~)I�>h�pAfO#�0]��7K"��x�����s�0�	1�]��.9��X�j�?�{o��XXƸ��tNp���wk��PR�"���xR*�6��\��a����J����s#��5�ĉ�q��!Vyq�����ξ���Uѻv(�~��#�kZ�_�0���BH�5	Y<���ェlY޻�9�<:������W�3c��S�8P!jQ�@l!�.֓��g-�Q+"�E]�9����z5f�	�|7�M�!p�lU�r=t�<�'1Ж�����^�� �b��ӂ\Ey��lBqm~�DD.�V���62�6���5-��t��m���6�j髎����qԓ���!8��aĺAm�{1���7�����m#�=�{��uY�R��}���37�T��.Ŋ�EY�|�k���zW�O9�7�d��'�9���#ƚ��wsR�KN��P������'e�ob�^����Z��L�bD�ϗ�'�h����xņy�u�m��SwJ��=/۫��X���]���}�0l�Q����j�` ��z�}L��,V�ܦ}���7B��9��d?���^�m�'gN��U��çŌC0��2By��Y+0�>��S�0L�0��|�����#�:W�n^��`S.�45��K�\Ea��#���5iUFw`��1�~W����)�^�y��Bk���@��v��7���2Y�l],���>gW��e-����6�Opf.LD&(�"����\���۰�6
:��d�|y��QH1[)��y-�4Toi}��;z��W���D�h"f�W�7�1��{`ŝ��+��$rd��R�Ν���&�--f'��{ 	�淃 7~q+>�
K�@��R~@�}FWE �@;�^�}{?P�<��,��uk���R9 �4�J3T��GkY8i�����J��(v��|l/P�H��Aٙ�q4s��_<�A`��)-���mo���0nU��'�f0Dl�b���K��_/�}�6��/�\C̻�1%{��E�dފ�g\8yR���!�t"&�o��Σ���;
��W�s�^IN��l#,MCA��Ք�Ƈ���av�&I㐙���%���\6�<��zP�\%Au��H�~�Z���ض�\��wxf3|K)j�������Ư_�g]O��AU����#'^�_VIv�J��;6�j���*#��9#Q��;s7+���S3���"���)�*DW�Ժ��
2�VNڍ��
B�^��!N</���G��稽����/�(c8H�~�T8;�^�-e�d͵�ma�2La�Z��j��q�ɼ·��Gޗ�h��j��]�4Q;{k�c�R�;Be|�z���V%U�$���T��Y���L��=�m�\�����󘷐2�~KR-�jF��XG�ќ���n�O�Gu�!Ԉ�ݭĐ _�79|��YM�HvX��,V�/�Q�!U�����+|��,�7��9�Y�zz�r�?�?d]<�]�ץO]J��Q�jJ�ޫ6U��-�>�V��.B횩I�֬��V3V�F��;�}�>��_�i�s_����s�+[	|�>�%�P3�%c�n<������P�0R_[����(L)
�����Qb}��:�{��6le���B�� jaq�W�r^�8�ҩ, V��9�>�}��_4Ҵ�Q0Ǩ�����/+?g�����2}���O��S2
��&.�؃���<Z��e�C�J�E.�_���Ư]��v�ƾ��d�Y����3�TŌW}��{o�l@�Qv����Ė%�0,�cnSY[���{+S<��\�j�K'�7�&�/�B�Z��/M�y�u4U����|����˴�j�ٙ0~\w�o�x�DR6̜v����7�P���F�D�6%7�����~�{� �� Y�"�MG|�4o��[a�̧��j=��Q|/^܂;�39c��2�8����vj�#p�C�p���:Q��Z��v�fA��[:s�����#!Uf��59���;��K�^-ާ,�T~��cH�s�M��-1�	��yy��EE��
�i>W,e�5��c��{��s�U�#-�j���DR$e���Q�@f3Z���uW�N�75�u�Uau����T�7n�.Q��\w�7�:���G���[�I�J��\ ؏��vx��* 2��*�]��F�2^ǮB����צ�.đ���*#Ȼ���:@�cjr���[}
�YџK,�m~t�7R��Ao�����p�b�%t��a��i�>�ٿ��x:��eo�L>�����)�n�.�ºE���o3r��z�<(8f��+���!�)`D#열}�B*8KUKy/��'�p�Dl���!�2��(rDZy�KP��ߢw.� ٱ�/�.\���;e���6J��A?���3�[P�n���>�V��s�N�M�����;J\�϶G��}�U9���z����)�l�T�=2���ݦ�'B0��(���W�ն�u��)��l��DY�
Kx�H$�f��������'A��j@ɞ!�g!?���S�? "�2GC��K+N/�����i*{{m#u��A#�&�T�ﺳ4��z����.���۩@=�}���٫v�"�fu_A�`�W�bH�4q�D�ee%d���4R3Z^�y0�}���Y���Ѱ�ls��|���nBf�Mt��~l\|F�)$�U�#a�T�i��9lj��A-�%���a5Z�K7KVe�XٝZI�ڃ3����	�%s����]g�*R�R<t���_���|����ͻ#�1���slg[��Õô�ή2G�f�߸T:z�����b�&k���[s�%��O��� ���x4Cx�}�׊
9-,@�m�h��މ�;ե�rQ�@�!-�������'�؅5�D�zJ��d��	3�����ݤZ3�sr��:\*UH��j����٥۸x��	"s[��4�㐜�;j�C��xE���t�S&���Z���c
�����N�H�b�JoiQUMIe��5�r�Na��bM�ްmɋ�dlx�k���:a&�/����AV��ꄬa�J����@��z.��$�E43MX��C^����g�:���F&Ч{�����̰���>��G#a��,�a?a��{=F,��ͷ���6C�Iᵞ�>���Q$��d���w�����5�q
- �Y�u�8�R��d��s�ܧ���m�@K����<��.����H>b�@��D3�3`h�Äa�er�v��)����y/�M���Z�e�x0L$��T��L��N��E��EH�oY�-F�$�A>�"zF�#B�~�`T�v��RH��>���xq�ؾ/��:�b�rqN��P��v�"��%�h_��"���Q���sP�+\�(�^�mXo�e�Ȣ�1S�U�W'�s�o7w�"��g�M:ǥ�8��$�����̼��+���];�1�顝��q|��[�����j����fs�-9.+_��TEr�WV�՛I�D��${5�?���לƗ���4�]����5��.��{5�gN2��fW$�IL��2����t����,t�x�kc���8��P�p٭�u�|d�<s`v���^������7�����j
W	���
I�E���233!ի�����~�ծ���\u�:��!�m�d��Y�f^Zؤ$�a�D���~O	4�'9ˣlUJ�A�h�,��6�K���k��k��K2���Kf��-�l�Ni��e�~Sm�jw��YV�F%t��v�}�� �'H��l���v�G�`��WHA�s���u���ĝ@Y��Y0�sW�h�N�+���WuW��'�����EOQ]n�]�=,̖��� �>QZ ���	tw�����F/�e#����\�0���ξZ!�`A��yƢ,)���D���C���6�9�P�[�K�﹁c�^��9���r��B�8h��P���\J�
�M*�>P��%a"���\I��۶��:^�:�Og���#e��P)4P¸�b��!�s|��\��ߋ����*�� ��ر���1�l�+����vvR3�f����߄Ev��m=�$��7�0z�b��&uB� �U����a�k0N�����m��D�1�!/�����OLH3]0�X�e�4=7�|A��L�t�~�4N��n�6����vO�7�"w��N��~nJ�4;ܱb�:Z��t�wz��# -���E&�r�ȯJ5p4P{���\+L�3�``��t���'����k>�.�
�Av��L_$���>�Ֆ$v������*܊�x\9;1�#Y8t���}+��o��s&�TwbK&,Ӂ�=��9�AȤ��� ���lh��L�kKM�b�3��V�ړ�ى�&߆v��h��GU.1�W>z5�(�u�l���}�"4W� ����AY�� ��[U�F�Cc���z���+�A0tj���A��?��O^@m��s�i ӻ��
���&|҂}�Z~X`_:\_k��.d���֫��Ѕ�>Sr��]���|+������Y�E�p�Ž�_!��ڬ������'}_v��o����n{{�Щ��~i��*H�'zVoŻ?�NU��B���Y�\��p:@%1y�1D3��4r7�r88~�OS|���|��%���x׮Y�yuB��a��/a�-����v'�ƺ�F�
�-��"-����P+c1V	8��s~�"�Rq0y\. |Tn�E�w��0��i�@��<7�$�)&�ΐZ��,��Ӆ>���L$�V�X�o�
� ���'ԗ�|y`Ǖ'Lٷ�r/@Fi���F4j��x"8+ʣ��Q�ٍ%��mI`�EC�c�>�e����I�$��L����mWKh��g��uJ�%0��*���/rV?�qQ
^��Y2�,{�/4�۩���k!!�q�]�}S��jՂ^}��H.��^���e��6Z2�F�Q��sն1}��ir=�i����� �����m܉A�>y`i��j��Տb�*�lchZ�b�R�Dw_+��<Ѡ��YYٹ��D]�	>br4Z��'8�K�����K�in�%u�Kom���E�b�b�5������
{���;�Zi����� +�����B�b�\�GgIJ�U��<cl�U0O�^�ɻB�W�=���O�Jۡ�z�K�y�=���Λ��V������쯟]�y� �9�InD���ҏ��]ow���3��c��/a|�GӰJ����=E2����|���Z�������Q��|}<m��~����f����}�u�����>�s�7��錾��g6�j �]RNW��i�-kLKc됗=��~QbcQ}v�LJ�
��}���1��E9��\��|����f�!S���;�hbAf��V���/.�ښ�ln�����6��������go�a2�^��_J:!��3���C��TAƅ:I�S��f��	i��eg��%��@�)�PJHΣ������5��R!Ͳoŉ���1����{��!�}Mf�9I��Y��G�����3/a���c`p�տH�x��_a�
��nI���W
w� XM�d�%̭����׭.J�j��r�utd�f�h9>��ܿ*	�f62H=wE_����f���Cj�Z�8w�a�)4�-��l���F�+k_�$U�2���D��8�X��Rߊ��ooFX�/��4�w�w%���I�r;�R8-{��.���m/ը��]w���=����b��-%�V*��C�#,�޺̳P���᳃���3O;tJ��Щa�J����݄���be�6���Z�}�B=�խ��̮�lOt�Ti]�zD�x��S�u�L�������_ުf[�̇c��N��5��F�$?�O����uw1���]u<<�(_��0�9d�v ^�,�rd��9��-�r�+W�=��9���!��!��rG���b�_[��Q��^�p_���ʂ�>*	"h*Mu�tX��+!\-�q�>L���0�pG�K^�7��זQE;�w��6��{O�&JriX��AB��η�L�
�1� >� @��E����vG2�O��b��C���8/�'���C�����,O��W�
��e�}��;�$n�<O9�:�g�!W\P�YW����'�8DErqju�]uUֽ �`r����)�+��Ƶ�AUz����)gz��c,�	Ԑ�1a>�Ý�v�QL%�ōH�� T�����`�z�~h0$K	 N��~7u��5yY�	���ާ]�5u�糞���nԝ��+Uba�l���\5R(��><Y�O]y�1J��y��J%�{���7��҂ǇX��	������|�ku���no���r"��m�����j��G���,A������k�l���	���N���.jՒ��Y����ݕ��7&@n~!�2���
����oy���w7��]Z����Z�� �>|֡��F~b�І�U< �&����0�_��ή���u��4��cU�W	��h֍����c�����&Lh���@��ʹ��Ud�]S0?��N4ӝW�f���w��"���zRl1�C^9�)��x�%}�ť6G�s�J�g��`��Uj�0.��k��xZ�V��R�2��4�$�Lᘊ�^�kQR��PB)4V%��F��Ck��[߾V.�Et%�#wO'������k��?Y*�3܈��Zc��{��ĳm����nH{[|)�E3�A.H�C�V��7����<�q먏
[��$���,���a�n6b������.�қ��(K��ͦ� ta���'��K �%e�I��
���|�r����j�P	����XG�hzJh�0%&�Z���S��~���������f��o������r9�ky���n�?��A扒҄�*����V�4>��4_'�5�A�4�ِ�� ��Gofg�6�W����og����Zn��T}}��7dgN�w{�����ɨ�\O��z,E}\�V�j�`����\�E�G�dI���.R��/8U�l��0�10u�K���&J����Q�����
����L~ڡ�{�����1V;����h"&v�ϨQp����o3q^�E�/�3�mJ�K��hSE���;	�%��O�{�9:x��-.��;T�m>�C��-F�2D�w�gl��&��d��L�­�(�_�|�>-�y�R� Aw�ǳ��K3��	�{?�B)���0��^���ڣcq]���9����O�ad���J���#w%,��biF-X�$�{�����V(�G�{��c�[�e|�(c�h�i�����`�䉽�^��R���CC]�c����+0���lF����.���w�)��Y�r����M��W��\��t�������A���01<��ʸvu�	6��^����u�����!���܈���Z��p�����qiX=���?8��9ꋚ��A��m�i�RZj ����	K�\O�CW�Ϛ����Ҍ���Y�=�T��_n��u�:�D�}��h��{�z,�-#���k�l�q��N�E�l�x�����ch�c����זcG빑LQ�%J�pͣ:����g�e[7�6��b:���lݸ��jh����z��gӠ��VX��SӚ^|��}`Pm�}�/mp����ba���=*�l̖ж65��o�C�_�G���B���U&�<)�L0�D�Z�2X�V0�w�	I��r=�c�&��=O�,��Tp�´|f�U{���l��pA3�*e�$�����3j躸����zp_��r0��Z�"����[���}������6N-p�z&<}�l�l�ӊ������-��u���^�����5Q�ꢶ�/kl�?�'d��-��M߲�{�YT,!kd�>7m��8�簇���(�q�2
H?���K���Ǜ���*g7ܭ���=?�X���̾��i������#��( ���*b۪K�'5��6o���>av�i�V��ѫ>���-���9�O ���|�f��z�;�/b�o���2>ћd$�XI<�(���R�pa"�	�1��|�Q�"՟�Y�}ݬj�R�#�(��t��!b�/�m&��vt����t3�!7_Ys��P���<iAY��G�VV����X���-�v���Ძ�;n����¶3�������_�M��d3iY~:�됐��2�=�Y�=U����L�q�"��:���~�i���OW�;�2A��+�}ms)׽f��]~��	�N ��"&W�Ր�{.�w�2":������st����y%�.q��Ϯ	y4J~$�%�� X�νR@�L���Y���+:P��-P_�~=���!`v�vvffx��%��{cQ	�yZ}n��&tg/�g�m�VZV�C���7��<ƅܖ/="B ����\3X$�mDE��77�-��Vwm�� z���g=���\X�'\\��NNb��T֗W�)�3��N��������1G�S]�Eo�!,���`�վ�V����_�b��1��������� �=�25~if�<8~�K˴ۓ�Vt�o�[�_� xX|��j�]ʈ��o�����^(e[��s�ſ�Ϭq�f�eh��뫪�j�+�aԟ:�zy��g���W��p�:i$Bh�HL��w�����/-+ӂ�#M��u�y��]{�Zs����)�臰�tݣ��8�=Ge�ݬΨ� {T���p����(�7�3��Q!�I�y׷l��ց	�4Q�h��e@��Z���J�U����D����NZ ��/�hkk�Ə��q��z������~d�\c���ԙ4tm_�(k��X�nC�9����[տ[��5���h&��C��v�	]�gOނ���2wׯ��s��ťO�K@m_��k/������H�`ڬ���#�G� �H������okC��z֙s'}v�
�����R��#FН�1QQ�nb��m�R�ʴKn��;�%�F��9�b��ΦQ��l:���� "���X�1Ħ�Fs�I��OdDE/iww:��TPv�y����Xp��"^�% �wo����U@���Yt-yv��3z� p>D��z]�] T��x�|K��/�S�N��O��4q�w����?q��*
�o{�,���s����!0�� E�s�\b�ꅘI�+�������z:X��H��I2�䎅�*�4l��Ď�^:Z��a�b��A=L>P��V�s
�w7�NLu���˯���+����V���&����[K"�f��VB�����XT�輻��e�Mx��Q+Ú���|U��fa�S�5�rȗ4X�u|l�=�=6���/u�3��X�-t�4��z� {��?�У��G���@�(-�4�]��/+3zf=K�#��y�E�W�qY|Q��#�E�zidܘ�",��7�}t�0�����Ҳʝ��.�o���j��Y���V�E�"�8k�/�H�2��]E^޸{�!��Q�DVQq�[+{b�J}}q�� v�$Sj�bY����:/9�ܑ�)�_|�<�����j�����b�����a����f�@w��g��מ�\~��:�E�'�_��iƎ�0��[|�­/c���'��f��\P�2��[��P5�`���u.�K�G�9$j�us[�B��W�)���O�������~ m��C6�\^a�[xH�P[lKFf��� ����
����=A����D��E�O���]y�X�>�����ь�/�mh`y��j��}�B��ъ�j]X����Bj��[x��1��.:����!���EM�-�ϟ}�Ļ�G`V� ʹ���5����av���7�ӥ���"� ��l�4�A���;
=B�5~���f��s�!+;�/0UaM���� K� �z�o�
,�Z'2�&�l,�x�h[�_l�:����N������L�~ݶ�ԀVzf�\�&��&�����%�ϝ��W�Z@̌ra�����K3�`�K\G�Y������M0�͖�I�i�~�tq!���3͝F�ڟy���tYt�����f�;��ɫ�n��Ѥ���-��#�F�4�)"ne��Fk
�N>4ۼ��J����P?dq��45�����,�0��7]q`߿���}�*2" .�N�)6ZK۫#��2 D�ֽ6��T8��c!b?��vA
���3q��^���V�]�;�m�ɽn��o�Çu#3g���ഭ�~�'πH���j��.�y@�(�я:���e.D@�%n��z��Ƭ�bGo�EK�XD�@��S*иD��Íί/d1`2Q?�]��*d .��
�!�U��]�t�Q}F��z�V��#M�ҵzKڲ�|�q�s�RT���z�s�-��c�
��!+5��p_�V�ݺ9��O>�����>Ar=�Fs^ Ԯ9Q���Y� 9e��z���E6�|�zn͟�}��/+z0i�,�|
OSA�!&�p��I��#qs���LzE���e��˃}�����1��HpT�`�0� ��$
6{�Z��ʫ\]O]�b��*�O�YW��$������R ����[�{�}c��J3�;�X��J*��mg�$ _��Ԕ�u�p����a��xT[�:���N��LΚ�z���[�9�n.�[�F���Z6�Y�j��ou>c�&��u��	���6��P++�Zoo���^~|���;$F��� ��v�y*����/ץ��#/�E@�H��Oʲ�Z�����M�t�-^q敠��R�!�aOñ1Sz���p���0[e[��V���:�T��?i��s(�)"�����_?w�l5��b�CY�.��œմ�љ�v�#�o�Bl�̑yke�4Z�}��rW$9��m�Mm%����pr_�Ď^���dD�h)� �Ж-N�;�'F߸|�>v'���G�*8������[e��!��@Yx���/��=b�>eAW��Z	$P����ܑ�'�w!�X��2�b���I�?�t� ��]�K��	P��\?'���:��WB�r�r�`����a���a��gT
����?���B@���?��70���`J��?B& H��k���=�n�\-�PP��:S����^��Z����{lr�8��s|��Jet]X� ���@��$_�@�ܛ�7��ׇ��B�{`.n�e���ڕ�~/�Ie9y��+g�V����rSM��2/�5�lV2fm��Wx�~�^����
�U��e����
(�%u���g�{@�cE\^��:�"q��:c;s|ɓ�I]'��x�.�N�����4�\wj�P�icC���70��@�ў��A���*�]Ө���l˪����e�Y��ʎ���$K�w��P�\d�vJ� (����Qb4��g�q�^굲LkfS�y�'e�,�ѻ��ۯ���"���KB4���Y���#?<]�������� ^Pie��ͦ���M��P	H{|��_f��4�?gFW�^Df���0�oV�����ƩmgS�L���ײ��^�S�	��Ƿ��훿r+��uX���W��W�ׯ̰>�Hh���AP��D��2[���ۡ��}��z$�>��D�#�Gߓ�:�jd��(p��^�̖=|b�8ю>��^��RR�^��4'/�iΰ�E%�E�2���pzD��	԰O��o��h�H�J��f�TT<���٩N��4ό��l;�'���M�v����uh}�V/0��ݏ�85_05,���XFW.�i#��8U��e�z���֘�l��,*U=�څl�$�9-�{A%Ϳ�@�� Ƅ�2�����Ig�W�I�3r���r�Y���{f�/�>�[Wx
*�_�P����T_���/]��l�R�m2��� �h��������;R�����2�bkS��4�=����)��Od9������ J��w���&}��a�@(�l�-� Aw^�۞���$�Pc�V9���+{�O4Ocp]�S���¡����=�k���Va�WyC�ʵC�p�)���Q�����{��D� �K֮���DB����6�g����پ�T�!!�a�hsII���/**�w�>)&@�R5ӭeǩ��K�?��%�Z�;��FT�-��� F��x����륂��ź@{dt��z�`�	��{4�[��6F�,	���@
\���P?��'��y�*�%�@�۷0,�Z �P��X'@�C_K]�������~R��TGs�5zDnv�G��*�˙YY����͉B�D�|���SQ=p��62r�}k<fn�{������� ע��A�N{�h0VU���z����Q�_��JӴ-�ݕ~�ڶ�d8o�<1�g���<��������yc�M>��Z�ǥm���~nJ��r<:x���Rw�OG׸{��u���@��Ľ�k��F�E�ϳK܈T����Iq2Я�t�+� o>���'|�U��؋F�	��_��~�2��I�[Mx݀  �/�Z~�8��[�.���c<(�*�a��tI,�O�!�d�f���R��پ� �	��aH{"H�ѻ����C<~nG���E��0HܷY�?�� >��������1�kg�+����\!��r����#,F9����/
Pғ�(1 |u�!�	���_��hN�V<����Tr� B�����%٦�QoVN?�BV��6��N�<ÌT�1~�h�f����b%s��>E"d{�cF��aW���Xn~~�����,��xl��I"��8��*b�Jz?������s����4�b��2��o��I��P��o�j'k��[rWd�Bj`C����+J�×�+�à�-d��֛���F<�:��s[SU��c4T�K<�r��!�W[j�=����?�<Z!?a�~�7����j��\/��ւ��=7B9f	��!|�'-�����_�YM�/�C>�_+>��C�f���V��'���G�@׼ ����|��5TTy�0���e���r؊���13p�#������>7�)��ZfA���x�94)ˊ�+KKl�_ߣ��ꇝ����G�0���H&_mj�A8y�|�L2,���EY�	� ��u���>�%"M^���}�H���<�Ѩrg3�d�r?������^�jjX�2nV+��m��&'�E�6,>�VSS�FD��SeRY�}�;�5�s�b�~��xF���r��4M�+���v��� *Ŵ⋚1�`�VR�^�Pv���w�g��ZNN~�1�^,)��C�J���܏K@j��K.:	G��ƥ/�A��|���$�6U2M�fj�h��X��9�������q��	@W
{<k��,4y��ɺ]��p ��M!��A,Y3;�.v��0�V�L��=�O/V���Ҝ�ux�(���AH��^�a�r�/@/�`ԇS}����~��}�5Kfm,��6�g����a!���[zs��QJI3���E�2$��7�˵��m"W�ʯ������>$ܑg�f�#y;�鍊�)?�`��n�B������!�NZa9�S/�P��2��m����[���J�҄1��ƺ=Py���sqe��'�r�������igg����W�9�;,���c�2�����S~� ���2��)���F��8V�^n�#��>я��c��P	�!�(�6e�g</<]�)�!h/���#�J�l�XA)C�Z�ur��Cc�)�����wr��O�j����b)l��vq7|����` @r`�8`����d߿��4&+�D�>�t�b�(%�^�\p?E�����B��L�=��^���"�x��_�_g&k�|
A���q�@3�S4�+��>ђ�^��͟�Ǵa&(�8��`,M�4��]�M6Z��M˒f��Q�׬ *�����!��b3ٮ�>���9�BY�,�A�А�k^�t�5�uie垴ژ�a�,���ܾ��J��5hB �s[O���##ξ�xxy��s�1��*̈�!�P(��WeF����l�����s�埥1�+�g�h��N�.�G�ʟ�h{���ˏ�x�}�s�}�Y�,o�ׂ	)v$���Sg�HW�E�����Ƙ؝3���/���b�S�}�N��=	����d���3���b��>����������*�׀�8qB����5�m��'�Ā�%�5Η���Ǫ#Yx�Y|)\aH̚�'���M��z�o�ψ��Q-�9��C��_X��?D�-�YdC�me'���A٢�y��
L���IS�lQ�E����mX�(�=��J+J�DT��S�Φ��1����ѽ� ��$�AC������;I�^>�3pǧ��ک��
�F�β�!;"�1�|���|,mXXH�*f�����4�;����y�O7�˪ �	i+U��6��`��B�nKĦ	�bO���4�<��mIg����NۆW��F��b�l�5�Ļ/��X��U>��B��A�C9>f[N��RxWgcv���ϡ��B���l�3������zX~�;��}�z��h����2\�rǉ&�4��hy��y� ��ZCc�nGzJ�EhޠC�
ISO7��Z�9��^���E��}�؝"[$t��tuQnceў���%@��.wBh�������w~Կ�!,rn}=Z�K���ȼa�3��������	��^_�񮂴��:~���q`�y�������X�A#{�+��@��d�QN�]��!R�#�3%��B���.���&׊WQڱ�T��P��n��kF�km	�N��U��ּj~R�?r�s�s[��n��Q	>=ڬ=�i�
 ,��dA�c���>L���,�т�^u.�~qcXz��ٽ� �1�Q��o��\ZR��v �@�a���7=�r;%Ti� =������}�/��6�\����!�7�Ty���y�x_�۷�W���f�q@YTV X%�= ���~CC0��0ɂ;�§G��K�!�p�`��ǻ�/z���"L��	ِv[�oO�T^�S�e�J�0
WZ�Dppw�k��<`ra�]1�&u��#/؀���;IqR.��N�h�s!M�}W,�3�s_���8:��i������dc�H��~�g�4��|�rO���|�/Z8#�xף��S5��>�
x�ȍ�C^�� ?M^>ޜ�����#�nU?�o�*�s���q(e���RAH����~>5��8���d(x��#�M8�Kr�4`5^,�{��Ǫ9�Ƒ�9������~\�S�h�x$.Q�3
�����抴w)�i×��U̾�f��;P,�����{�J�Ң��e,�,c?7�3��L�8X��p��-�3���[0����zǵ�� "�-52r�~�ަ
we�ߎ�����X�jR�tHhQ�`��uE��-Ь��j˳�T�>@a��N ��[�y��~��Z�큥Eqή�T���[�ߛ���&�]xܻ�.�y��Pd�Q��M�@ ��f�\����{�mb��R\�ב��ư{���*�EJ�C�cr ��C�����P@�
3P�:w����+:�٧�핦��BS	u%ɏ3R�rн�Dt�\�Ƨ���-������?n�ɿ��^H��R�|�C�m\.��~k�#���𫒣(3�;e��K�Z���_�hP���hO ��u�m�5����'�bZ�x?�Q]W�~�@	��A�ƍ\�ie�.J�hp�2Y����{�}��.E���3��b������v����t�k�5��;�#�����c��u<A�	M���֍Y��t�m5R�_�WG���[�W��� ��izy�}�z����I?p<#�E�x����\Ϊ.#9�hR���E�N��wO�c��ݷ�^�Xٽ� ��JT5���zPe�C������ �*~�_u�a��j�(c�$0���Ё�vYZFܜ���2�e��S�wGJ����v7 ڻQ�+v�3�!��	 ��+s��fG�����zX{��_zɈ�s���P%#�:켚�^6�]v?����ȣ���g`������|����>�!O3�g�Aa>���Ϯ��D{�y�W��T�^�\�B\)6�@�k}�#�	p���_3��׫i�|RN��
mge������10��BVg9��i��W�d�����GY������ܽ�r��m���r@�
�����2_ �w��L�?��D��;�u6�6���p Q���R2�&�,~K��,L��&6l-�[(����RCi�H�ce��*�x-�T�e�n�]:�+� �B��I��R�����9�pn���$7�zKXv�&b��cKs�#����|z��%�9�����V���l
�9)9y���Hn /4b�G9���<6Q*�q�k�1[2뗛�}��}��#��bE�\�p�/5�DkGb*�Gpm �^���{�xYQ`DV���F>l���.���;{R��ĥ#|�R3<L��A���r�){`�����u�>**���+�[*#�W��^�dԵќ��j~�;�K�&�3�+�	���ЎciV]��	㔘��|��R-]��NH��y�U��	��G�K�#ǄCN�8�X9c,gI|}c��xP�'Ι����čsj�C�m2݋�H!���
K�e$����]7���h�������MpKW�9���V}���%��$��&����W��~2N��}[�e/?{���ř���#��/z��h��K������00��F[��d���N���D����>��]�]�;M|�O����d5�����:�`WW�ǲև��+9�vt���5���q���/��|�l\aP��#�q��Y���CGv��k�H�	�����!S�\G�Z�^�K�f'�;NW<�T��.�m�2|�7��qLA���xEV�h.qC�b��v.��w%��=�6_`�5��S�`o�����m��o���,z�O�O�GZ�\]a��xO�c襂K�#;�u/[)�ǆ�?�^0W����H��ɿ����Y+M܏����N,�@oT�{������E�P�٦�oP�7����J��@�Á���@����g�����gu'vC��g[�/���/�&�^�/��ca���Kњ=V!
A01���K>��褨��k�� ���w���Q ��Lu�T$��3LO�*��Ժ^�)W�yu|p����F�AQ񆨨>X��O�ϟW����x���1�/Uv68x�5}j������
g��7�|6/<HA;�V�l�a�����s'xA��Tt`�l7"9�O_ �������dL��zf�>��B�)��>�܍#�$~}��c�ac~-a��q^|�>���NQ�d���v�� �G��G��5H/�T�:r�<��6�߶ď��~�K慏�3�DO_x��a9�<d%�#g��n�F=�z�������'�Q�
K�m���s����?s��;˽Χ�q1���Ik���k��Zh�S&�uq�P��\�����(	��hgI�m��D�q3>~���Q����O�H�~.
��� +���җ�����&��4a�盁�>r"Ë'������i��KAf���S�o�J�!Ⱥ��3ɜ����(Ǒ�k/�#�w����#����	dQz=�+s�|����xa\L��ZĜc�N��`Pj������s��6RQ��#2k1�]n߸�zf�rP���Q��eXX܂u��C��� �z��$�X���ɤ��W���΄ג!zNS���E���K���ш���ݎ$�|��]��n�ŷ�Q��e�u𷺩Gޯr�4R��J���ڼg���-z�G�}(lz���1��K��yu,�uA�l�c�H��]H����ޙ�m�����/>[��v��K~-����K�#o`�;�x��sE�A������� �K�*ɤ���R>�o�9=�-���";�x$��D����ż��ok�L{R���d�˝eە�� ���p}qTe��5_����/�i��V�#*"tq >ܑh�ʩ�zQ��7��}S�������|)8b�OxiM]��K{<"j�1׻��T~ʒ����5�v�߯_�6������Fms���R��}Kv����:=�N�"�g���ǝVO"�f��	�%#��`40�\���i��&Yp#[���%����D�{��O�f��;'��}�NlG�ov�=�[�C���,*,��wi���!T~����{��Y�Q��OF{w�"�N���}Y��i'��t�����E�a���s�gu/��c�E�T���_��+��m�ii�<p��_Q��3ѿ'��]\+_,����4x�|!C���č`�!{C�M�>�˳���/�Gf�ě�b.��k	tJ)rZ/��1�&}��U�Q;�g7V�$��a'{�帯qx�Wrf�I�Z����=�<��YD�G`H��/w�x$��7b/�kj��/��y����(��=���3�?��7#��,M�\���`�gv;�ZC��~��AkZ�N������-h:!�-��E����0䒲'e|�cHf_����p�us�f!����*z{���z9�/���e"�̻MϨ+�IW���ҭ �����C�T��0���Z~+�g[
�H�5��!,r4��}bvG���SbE���F��ҧ�g��J�b��q��=>�F�,�
+�^�V�;}��K}׍����}� 8t8�n���4-�a�R~Cip��z� ��fC-�1�rq�r�
 �=[��r�����]Sb>�(It;�4���x�)��XU�O�{�=S�B"��;ߞn^F��F3�w;A��:rAN��~�$ێ����h�75��p��O��&?=��;�bk;�J=���i��EEV@�0�챯/�P��R��C
�7�X%��F�Ip@����*X������� k�m�x%�WAr��` �#TD���K6,P�����1F)��I�6B:6�e#�����}���C�G��㺯����� By�2���XW�N(^n�!��6w����*b�3B}�@��=���֣��'��6��]LaS'��Rl^����%���1Ύ�G��[����[SL�­i��	��1��@�E9�s+s̆�5��)�q N��Q+��<�ō���$<>�e7�t���'�]�e)b2[�e=�}��(���`��K���iˀ�6���w"n7!}�,�1�mR���.<HG�)ud��$/�n��G�a�h�?B�;q0#�)�d��)�+��a�3�����LW3��oW6��?w�DL�����/��kO��A�������4�J�^�t�8�߹��G"�����ﾥ$��2���3|�7�\����cz���-��(P�DY����nIa2B���X9���Bia`� �~�g)��Z�����������&Q���^��O�	1�T�,�"`5����ս�T�JF�G���m�4�J��XC"CT���y��b@���i��즄"�@���Ϋ�S�H;x<א�I-�����c���Z'�
���F�c��t�)�z׻F���v��6S3��$�4�++H��bNe@�����{���DpD�����3 o�/���$;����7q�n��6�
����`�^T��߰��gJyU�M�49�a�h(��$� ?Bo��g�������"�P��`ݣ��K��wV&��#Xv�~�x������r�g=8���L�3�C�5���G��]�R)^c�
E>�+I�M&>�v��������e��<>����ʎ���/�P2
?����}ooѯY1�"tM�5�舫��$���7"]E�/�����%fVɔ�OA���V������ 07W��lX1��nK]�G��XM�z���/Pn�)~ۯ�4�)��w��b�|{�7.��1��⡟_lj)��a�tӎ���V�Y ލ������p,ǁ?<I�rE��֏�]��q�R邵3�Wp��E���8,�ʶK��m�X�H�<���'�xP ����V�@q�_B��?�po�g����F�"xi�&_�hƚ�h��$	�7��՝��ˇ�,یU�#�9ǆ��`��K�WV�]�z���_��g����%�'Z_����?w���m#�7d!C4���4����+��Ɔ�r��.���%E�j�s�x��	# ��q&MS/
Vz��a&���8*@2j3Q�	Մ�� g��,�OA�Iq��K?��֫q��j���>���I�|'Q�Rg�}>$���!��$��<7�PZN�@y�^����q	g����h���)KA�N��3�Xc6��k��Lܪ%�x�(�N:���s7g���&S���pT��nW�������V._�C��:W�aU�X6�~�v*��x7:R�`�[�����g􅂂��d%`�^7hQM��=i�;�R��W�0�ښ�B��Ǳ�w����\��Y!�D%��ɸ#{��GUb\2��M�/-���k�_-���6�Oÿr���}	Q��
�FH��2�����"x�A��;��٨j�
&!y_��{���\�K�<	M�����}$�q&�
u	��Udm���ZV�e_�P����ѼH/i���6dR�019���Z!��{7��8��L���'rd|����隷^�������&��s� 9?�TUA�e4���Ň���W�5"�������7�()���A�*4(U�8�n��SD�MQ|���& �s����E����J	�H \����ѧ'��rD�ʝ���Pk���������^����%�	�^��1v�r��k�7x���}(�!�R�
b�k�}c�g�S��sF��Z�nwk iY�DyF��N�I�F9�P���6}2$fK��a��Nw���e)�$=�p��Y�i�LC�}/����������%����(F}F>`�H�i-~H��z�'�����Ӧ��������q @I�!?}B����-�ɫ6�L�ɺ��1������Ke�K�����TA��'w .^�8J�<J���%O��� �<����%�TdK�V�'��]�¶4�=F�3W�|�W����!�{��8�)���o	�q�d��`�1B�y��鮊&���cYp�Zd�w%C�V��O$);�ݳ��߱����$��m5�R� ��e#��D�n�y�SZ+��U�.���a����#�[ko|M['m	�-�i�X��')To�I�����LLnR����n0��W[�������H���0�+8<�V�A�(}z��) ���gķ/�ø��#�30�l�?�뱇9��߻�h��Y�[�ؗ�1t�r|W%�����y1Ѓ6&��I:�+9�c��Tpݖ"���>D�;��v�%�c�1���w�Lup6W���W=E2CZB޽����a�6���s�Ҩ�ی�h�F�"�K��]��e��d������J~�����U�2T{��Y	�7}�?H��V6�!o���/��*�Z��)��ؚ���fU�h�+��y��g�D�����M۾���X���t���������;�!a#���M�����N?�e�PMc�K�_[�Yg���J�Q|ս߭�|~@5}���O��Z�
6&�r���M��<}�L��}
;��1�S��������d�g�v�؇=,6U�Q�U�I�.c� '��`K�CS!b��,*E�T�wߛ~)���  �}�}ݶͮ�F__}g'�1#�-x߳⧊���e��5s����^L�K��+�Y�~T��3�JhBP^u��������q�Ow���q�',m? �:�\]�{=AH�*T
��C:Ǒ��'��i@(�ԛ0�B0cL��~���1�N��\�s�|L<7Z�;�2�X0h$\��\�8 )�0�Y��r�aC���Ab�μ9�H���+��-r���F%�Q߬�E���E�['�#W����KoS���������{׎��u�VĨ��bo5X���I�%�޷7!H����An��%%�� n�����hRs���z�	�h�5M��NV}��ػ5�ޱ�6��,v���*��g���FΉ��'K��~��t��Z�X�ct�PW-*���6��i����ί��-����b�⤄��҆�>��N@�� �a,0d�߇a#�����ـ�i�z�y坤�����U�c�v#�^Q���]v�$"��BO[���R�G{*��r�N���+"w3�ݗI&{ch��Y�%u�UB_h^��ܴ����Ir:�o�~�;Z��ٙG5�N|�c!�n�[����"-m�8�57??���QKL<m����KUU\t�W��R�_�K�_�Z��^x���Da��g*����{�j�(d�1N�~��i����I/��];rFi/�֮�#�;^%0b60U�Bb?�QA���?P������pH��6A��^�ʳL�F��|�}�3��dB��2��T��A�vP9������C���sc�
�����)&�oD{i�7#=*t���p'�4�O3�	�!V�f�hc���p��Ya!��:Ɔ����5���D�!��ح��$t��R_]�,���z&&%����y
^�n*�����25����]GҶ.p�����uH;��^vk�e-�,+���3W���:���0��r�N�
�U��9-�2�#���7M�ބj��@��t�S��{���󾈺��Ғ�Tf-��w�!�A ���C���~�,��
並��8<%f}!�gg�]�튲kx�^�rN�J��]���5�����rWY�W��4v�,<�A�r#8'�'r�E�x�w5���Jh�[���rƁ��^��w����^B$;�-��M��3ѣ����2M����HX�y��vG�B�����Ft)���&���zӵUA�$�F�U����%���T/s3C	�����=qh�~����'��j�=8�M�SM)���6�_\ ��e<�w^��}������K�i�܌�C7����^���c����
���Y
Od�0OVo ʠ��-~��-K�D�j�����YG���f7
Z���kAȁ�VPLL����EFzH}�TwOO-����]�I�;�s��&A�n$VQ\�3���\u���q�y�A����,i�)�H����9��������)�n�'�@N�}�y�����d�'�㼥��)���ԍ�3ΖS*r�ޟ?߀���j�=����n�tgU#%�v��~�}�d�~�&��u6����fn�9��?W��l�c��c7��bUؤ�5>��<�U��\�΃�}|�����J@O?�:r���Z�Ĭ,�.s++���$��UK�t��i{�~���8~Ἀ�:(�*��<�`$�\��y��X�*�f�]C�#��_S�ݸ�?��
�����X��j����<U����j�H��g����D(g��4h-H��²"l�����i?�`�I�0����t{��{�Oߧ� �'���Z%
Iu0�9S�1ۚ���4wؑ\�p-����{����O���T�u>�����v��{p��1z�E�/X���n?�Jx:>f�ʶLv��tR%k(�6��������u� ]��J���YU�dJ�{�����)oX�+�y�R�{�r���C��H8�uP���qc�?!l��� ���#p��x:�яE�(���ے����;�Y�������}K{����Y�U� �G�C��zwd�,_�Gn<ζ@�̟�����"v�?�&q�8
�<sd�q�ȡ��,��l�E&婫.v�y�q}���=ZSF�:w�;)gT��Rtqj6��1,mSݨ�K�z�֐�<��Y���S2�lۿz���J���vq)���ӿ������nćO�Y�B�zQ��G2)F�k�?�3�Xq��o��z��ˁNo`� ��=������_�n��Hm�Jj�u�S�o���$�٦Ѓ\���Ϟ �	��x�+8��OM䨣�}c��g�K֝�FQr��ԧr�!��!��!�WY*V��K�}��(g��[c}M��Pi���$o|�9'���}�#4��.�ɕ5��Q\\�7��q�&�$Z5i-�COs>��gwl!wF0IF�#�?]�?��M�[���V�r䫏����y�[M#{�����W��==E���L�y~:��F�<��8ؐ��Z�M�Ǿ�@����4�uo�21�����;� �G�ZLN���^y`�@(]�?�r�v/��Vk7�����>,܏<>��w�N^%'�n*�E�5�,�~�%P�K%����y*M��q�HF!��yC�d�\�׳7���C�n\q\/T��Y�]���,
�����O%uT�%5x7-�'$2lx�Ll�<�G�%�u�Kڄ_
^-��ه=��D��ڸ�\7LK��&F��qXϮ�ϝ%��OXT��\�k��(�a��\�Z�'�O5u+}��O#V�,�wăy���ے�*OO��M��0���x�l�΍��L�x��D�))	�hr��;�O��Vϵ�&�DPpP�j�ϸ�y?Y��I�X�α���ޕYlH?rmg K�"C���N�'5���(D�~z2Y���{��ꈍ#�{�i&��tL�mU�Z��=���%��
�_Z�����]k���fi��|������7���o���}y�������A*� s33݀�E&փ'��Yf��Jn����A��)N����$ �Kh�w:���Iɒ�W-�ʟo��v�|<���B6u�|��5vȏ�?k�+Դ��<�8{���wq�,�S �^��mo*�y�<-崠�ù!qX�vA&3ٔ(���Y;�ʢ�@�:"��2z�����%�Ac+��r6PF$a�5��78����e��HQ���#����S1�G�L�[Lt�s�뙨����6�WkbK؏����7�O����:���q���~F�Q?���4O�n�Y���o)�%ro~�&���W���%�^}M(KrR��Rr�'�ǵF��Ě-ĖRYí�g�jcq@����HĐ_������ʓ�ݨ��OVA��zl���v/E+J?+x����>�i�	�O������Lo�Cd<�_���o��P�Wh>2���_�i�O!�h�Ĕ�^�5g�j�K�/����2¸�	�]�u�A��O�,��1��`���#fha�ԄJ�]HD�o#t�ʢ"�>L
�آ��s��_��;]���l4�B>��6�������>�����im�ݴ��ڐ.S��+�e�,?��ȉs/�,Q\�in��%F6��C"�do#���pD-�m<�^���xZ������u�X9]���]�i����12��'��m»����ǥ(	Wlȴ����3���fE��C]`{0�ښ���d��t�6yL`7R�����!���Y{{Tm��Cۈ��N�ˤ��������#�*k��{�DS��64�8�{��ci��Y٢� nG�b�j�M�s��_?S�u�3@NbߚA�¼<f��w<?Ň���k��nG�^���7y��)���Z.�gt�w�8}� '4k:�o� >I�X "����t���$#��ˮ�뻵,�Gn�օ|zv͎�'FWE8]�M�L8�Ze��� �W���]}�Q퓷��;���ˬ�q�K�o�^��UIg��y��6������{�c2i)����d��UO�W��>�M)O
�	K�R�7��#m�����v,�|�^' �g8$rO�6��G�LN��~������ʳivKn��8:�쌓�͒X:��P�m@Ȍ���t�^/����h�"���U�ۊ����x���w*8�k��^/���dxDM)�R�e�^��Gd����� �w����$��Q3��-W1uTɦt�B���OW3����Ip�0�����,k�F� ���.
W��+�P�Ҋ�����Ӆ�Z�"����:��;����x|���!�Q%�I@�쏉i��^J��6��՚����DbNpK��fL���wb'΄-��qE��03 �3z��׭s��C�lH���V��ո`:���Ԁ	F��4L�����['^��&����.4ASJ��=�Kj�ޓ��-R{p���}S��0�]
�<~�����+�
�J�3?x�RT�IM�qK��+*h6{��Ic;T��1��L�Z�/�o�*��뷹��q�Ir�~�� ݦ�(�I�t� 1�n[XeHE�������К�L��[ǧ�4o�Ŏ�RO ��Y���[#����Lj?�Z�J<|�q���$(�d�u'�}���Hͅ��ۼ=8O���y|�Hy��3^���|�/�\�׻qorIh��	��6u0L�^��7���Z�8����&o0�r��\ �����Y.22>tMnȇ�5�/�b-//O�ژ㋎�6�'�
��O��@�qӅ����y��AҏOU]
M&)�l��&g�R��5�GF�IE��x��>�;��:��}m���ZH����QO�J�ٯ��uC���w��V�;���K �eY�(ӓ�鸮U9=�Ն,w��z-�|��qmt*I�fh6��.���G9Հr:���6&`@��?�Ru.�VXS���N�ohd��.� ���A9wdcdo����͑L��65�(�6�=�~��ݣ���݊mI�Z�(��V�wU�ůٿ�h[�F����Nɧ��й�g���x��)|�|����Eq���B���Hzk�-���^n	��G	��cF��>���]�}���?�x�<Ϲ�t�X����T�n>E��,��M�����z�����m�@��;�����t�n�����U�W�\�L��'�c���rnqG?�z3%N,Rx�!� Z��T��{��\�������Gӣ��K��9�E��0�1̠�O?=jB��8Y����T��s��X��Լ�y�!�b�W5�Z����*.:�+H�k�K
�t������=K=v,K���Sw$P��tQ�b��_�]'�i�2���bw%��u��5������O)�^e��R��/���k��g�:o�4�?����W�e��',k� ̤�^.�z���A�s��{͡���cb��@�����pv�j��� ���HK�A��FJu�e����y�Ŗ�EXϟ����֦���	�j����	����$S�>�S3%L����Y�Lt�/�!e�+���I�#�jT��E��;)G�a�H���N�%�߽J��%����ҖnVw �:�O	;D+.�d7��r���a|��:#7Mk^�T5&�
~��.�e�RR"�kf3�������4��e$��@p�f1̺h��#=�ѱ1��]�5OxFo_��>�x�G�#�̎���[k�����ӧk�;n%6�7Q�ؔ~zy�|G���t0--.6�e�C�):5��m/͛7���? =���n>Ӎ;[����|�r�~!�*^V��iet
����ɕ7�s�ٺ<\��Ν�/�( K��m�I��8���C���.[퉫����z����S>��O♣7x1@�U���d�|�8w�"'�]�n=Fο���:J_���l�?_����V���y���-�g�y.��ֶ=�g���T!�=������p��̠��!��e����6�sӔ{��X�sa�L	V� ��-��o�TWT{;Q>-)+ӁB���au��z&�_�%�3�|��ߞ�*K���.���0����H�A�d|?#�� �}��^�/�i!�����e5d�&��ٻ���wr�"`��攺�[r`qx�0���g��r�e����q�#�/���?)>L�m �Q�n*e�ښ�Pc�p��*��*��~��6p���&�馣T'd��x�P���n��	B��|��`�5T�:�J�Z�*�V`%�TM�C���r�
��\����ᶶ+�Z4f7��sr�=�b��)����b�I�d�ڹ�I�]O��0/kN�|s��$$�]8�WZwJ�	���9ñ$_�>�^9ؕI~�Wzc!5��ʇfgS�6�������)����$-W��~΀ ۅ߆��諮G�0b6�&��::�O^՜��p�1�r��� Hd� �}0�Y^Z:�\�xdcj�������Wg�ϗ��/�prhxS�J�/p��:N���j ŋ�H�}v[����<���{E�y� �V`g��a_�E�:`�޲6�yr���x fUOxE�Q��k��x�;�c|�k��Z|`�����P]Aý���o!���b���&��%��>2.�t��n���d��.5��
��������;z���s��7gUWW�Q���KLT��yAm����+�NYj�c|���������Ru� ��v<`�Ge� �+nmQ�F�,[�œ�� �V��pX���o!���9�5�_ �t�^�%��qb���}��pd�k�FE�{�^H�>ae(��,��^F^�i���*j�6�Pn��S��.�j��2Ⱥ�b���]gl��jE�5Z'}u��H�Z�E�],wn�#J��B�)�u����^箾����S��������,5>%a8Xs�Ȱ�~�+����3�|Fr��.b#�"����r��O��Bwy	���eX���FV�:�d�n����SN�)n�<l��N��J�8"'KЯ��d�g�R d����'	��T�4�Vo:ĭ0�p5�ӹ��9۲164��i�V ]��M'T�,�{�_��j��m��P�,.}A���|��K��wS��C~���ҥ՞�;]�{�I��r�IIBeͺ��-���mj.�o�ZT4r=:A"��S� ]5E�s���۬WX^����T�/���Oή�������#�@�E���<Q\�J�����
e�Ci{�<">[{��v�U�!7��+�Q E���e�⨯�⪮�<��]	��D�]]%0��`��5�14�n{�lN8��Z��w�Ř/�nw�����w�����N�|r��a(�ZN���s�0�5ay��������l�X�r�h�KD{}���6�����sh � ��\д�����+��h-�5�VGΗo�z;k%
�>���ɺ:T�7�ous7W:��2��	��qFf4'������Ή�����ꋰ�a�Md� u�0bn|$���w�q�Y�^�<�3�P�s��M�&K���.�,�����|���G�2`� �V.O���In"��P�B��hʦg����rT����z�<��#��P���居2f>��gۧ\��Hƒ���.7rN�q�+��1peB(���?oZ�tlZ�h1۟��@��=l68�]�ܐy�.����G�,a7\���{�c��*6���>��8��=��m��8�;M|��	��5����8�08A���*��՝4���������r#̜A�
�.I}CQ��k�~O��b���ŽI�iw6��AǪq<KR�L�<��md��ێ����#B-��]�����H��N>ھ S�?.��nY�����Zaj	��j ��t�����O�F��=G�O*�+��Lz&�UȄnY�c�/�}�sn�p#���x��	I�;ޯh�U��6�ա�:��x)wa�������=/zjE��쉟 h��!�N���}��}5W��A�@4�VW]V;�G�] <�C����#����)1�zcF�'�L�)C�ď��	3�="*��f��=�c˿�m7y̲½�Ĝ����U�h5*�F1j��bڮ�R�KDT�8P�����y�XI�=F�ɪP��*�dU(��S�\�7�wrS���4�T�&�{ �����T��ͫE}�t�ru^e|R���������u��6[G1�=�C��������G�x)�	K���(���^���KP��٥�;�t��
��y7��0��vLS�0�mN��'��Wi!I�<�$)�������aq�ÏZ����o��NO�j���K�IY*I(��#��#���R���\V;�{��j��{δu�D�K�i��+�  [�(�@�Բ�Jk�G/:!�7SUw�S��5�o�q�+��7xSS����n��=BS#�l.\��8֮�>�F �w�&@d��r�]�]�N�F��������u�-����ᗂ�%.���Jj��颍��	Y���G��U*��S��H��'SŚ���z�4ick�F��o�4�3�n;�7��!h���Ti�՚J�<�PuQ����w�d|���c�6�^|ր�
�M�}n!'M�>Oy�8�!��x�h#�1���{���VY4#�*����0�<��j=8����8��ܚ�,��K��
��:r�g&�9�[���h����ul��02/b4_��Ҥ�H+����.#�f�DPR��[�c��Pߣ�$[c����Յc\��0F��j%����;�{2{�g����X��p\
�H�1O�l�O��ij��x�X ھy�"�4�\!n���Jַ��~�~"�+��&����?��Xߜ�H�$5��r���L�h"�T�D���￠ʳ#���>���GI�uu�%�����KǇ&f��R�3�	#�6r��8Q�#�-�RF��"[q�V� {�Jl�أU���mu�Ux���ug���R�{჉+��S	�z�;�0��b׺�~m-�)��>�>ʊi��O<�É�ށ�V�{L�(�u� 4�(��Li=��0_�Z�	%~�ى4W���>�[�Tx$��E��;�C[s��١�q1��e���N;�|cz�c,�M��&�7���Z�;�//�V���WU���'�Z6r�I4��l�Uc��[jc��ۛ����:����o��̑���}@�-�A tǶ`�fI-�9	���I�$G9�l<����U�  ��^Z|��5��m�O��O�9y��jd�Q�%M�!e����3����ؙG��>�(~1��k��ˮ."Z|^�Xn|��Jd]^�} �j	l��5w�@���gcz�BK�˜��<��;� ���)g~o��,Ex��,�!m��LΤ^+�� r8�q5�غ��,������v�L�����ܻZ�@�5�*%��@O-�=�~M�z3��:��^5o��6� �׾tWP�
Kזx�{�`j��s(4p'��^���+��<^�sأ����b�?��$��xH����zE�W�3�	J��%'��5[act������	n��hO��׵1M�0���a����M���&���:�R�υX:���iZ���
�rAM�
1��B��MJ�~���U��8�N��Ϳ�����a��.�l��"��_�,����|�t�N�h)pwG5 �^�w#4�3� ږ��=b�:� �g���*y�To��()�XE��PI��R�T���z>��O��5�w���|�ݙ<�ܕ�qk&'��˪m�%��Z*K�F�Uu}HV��@k������q�����w_�h��O���-�-�8�p%Y�EoñC���7c�c��w/�rЯE�m�0XN����ëؙ�x�K�ʔF�2�]Ru�f� A��n��׬ �ī����Gˉ�5�7,���6��~C���S���Oݣ���y&ʡ�Aڷ=4�'�K�$��)p�ր|���읭sd�������4�<���`|��s ��k[�da�ު4����7�t<�T�x�a %�[[b����	���$�Z�Ӏ��*� M���uGE2��ޡVTC̛\}:�����nO�x��ر�[�	\�00evBT/��az�����y���w��f�cJ�� ��?{X]�-y�r�!���%M$g]��ﯽ3Ps�����z����>l��陸/>:]�72�����J�+���k@fI[��\���&��~���UZ��� lle`h^X�+ޚd�+z��x�[��t�"� i�Q+����9yy�����@�z���uZ���!�aO�5&N���ڙ����Cӂ�bs���y�{�<��ᢳ�-%.:�7~a���"�����O7����Y<���������n��,+�!��x��;L2���1h�ȟ��>��[�����3"�y�����g�	ϙ�����?ݸN������Р�:#��&A����=?<��Q\�ʯY{F���h4P�B9	��?��#����_���pB�\�Tr(���L�G��bI@ǽ9�+��0�;���.���K�:��_��kB�q�ϣ�m�Q����������qx<q��C�T����v�߼�7H�s�G{�_���j�w2���X�_�?y��g
�/'��/����=&]^`2[�?K<fF�D������8�p��td���N����QE5O�z[�I}}�m�o�(��p���?}��
iCn1�����=~L.q�&�SvI��Y((����VE%W5G�t�.x#��{3F�S�p���d�(Z8�5���bi�=��.�v���&C���qr�(��L����5��ik<�
^1�oԂ�ü�'aeuV�!{/��M�B������͊�I*zp�н��A�+)Z6���Kn*{��}|��� �p�����ʕ8�?�����/����{ؓbS�����KZ*�������=�O�����J����{h��ڴ�j��~�����r��%����E�z�h7�Z��s����#>�qF
��^�@GCwM��_ۤ:��ŉ�J�C
�M�)���8�!`X��'�t��⩻G>Ļ-�ƻ8�>a�pV��y�o����x�[/b�+eǈuoĿ�ɓ'ێ���c�r3_��'u:���������$�h��.�+�o��6��R�x�Z��.��Ѣ
��A�~`�> �n�aI���Y�y��/+��)�#t�$4��p��xv��/�ģ>��﹈T�V��Lv�|V��~�);��������f}��?vK�0b\��f���͖u2���\�霢��p��&3��K��>��}��U�)��H����-M��x�2\f.�v0�/#��Auܠ���Fq��v�"�!��&['����Ś���]se!_��T��v�n)��#�;G�P�t�b+����9� H�q˦�Rݨ�qQhE��ɮ����LQ�H&7��i��ÿ^7���:Hˋ����Gna$�]0�5҅��#��$���A�-9F��C����\�n�K�I��0�.ov��zCf��;��p�߻�-�L�-��R>��Ɠ���Yk"Z_���<3� T�
N������� Ȳ�8e�Z�n��3�Vk�>\j3Z�ss���L�|�P��{�a��z��Y��5sm�K��UxV��:�x�;�ƍ�#�(�L�A�L救�dY9T�
Wi��NNQ����R��+mQ�e<^�/��'͕�wQW�C�uL�昿�|6��"�%��m�����щ�+{�����=Z�S�y��K� [�I�(�_���Y¼�G�%W�z�~�m�5W�^�$
�tgϛu0¥Yp����s�+�V����6*��V;�yF�Zw��:f���DՒ�6�a��η���4O���d������Tl���9�j����5�|$���!ܟ\~��+�oy�;b��󹝬A-��*���0bt��c��$�/���ӟ�b�=���b���������(vW�3%�l�$��.W,��"E��PO{1}V(��7p��חO T�D�_�j 능��~�I>���)3�<�������T�NP�J�� ��V����䥱ÊXڥ�7�&ź�v���3���y�c��w����1Ѳ�\�z�E�=

 �u���J��BlQ ^��(֣τ���E��])pO�0�-�I���g������Z����Wn\/�|��v����h��wrrz��߷�u�$���g��.�T�h�Y��g BIVy�\{}`T���,Vnl^>���v�
�]����;�X�#�M/[��s���F�:�mbϸݢ���A�k}i�����cv� ;�p�ۊ�^ʁM������L���&v,�+�DD>	���s]y� KA⏻�eEZ�c�hoXCl�2ncm����v��[O`��)�J��h+�u����6dgUV�f�������m��;Ɍ����P����L/�3F~��X�>`$1U���f&�@�����daޚj����+D��h ��9^R�2�bP�L����C��?{u�2@o�K<"{��JC"#ތ�>�>F=T�TQ���O)~-}��*HV�^�7Z����=�j���Y�rL�ܵ��a���_�4��,�k�2��8*�olq�n���s
a�������<���_���{�ӓ���|�"�9X����c�
,&�qJ��eĈ}�U�?$�	
2����U��,�ۃ����s�h��m��������8-t'��9�Isj0�S�./k98�D&����J<��!-�33+��74,���P]Ji@��cqf��5%k߸!^)jYh�&p��xA��*>���=�[y���������m�O�Y:�x�����u��Z�AEC��㆛
5z����X,'g���iYC��6b��Nzq �TQ�3�{�f��\�EP�W�	��à�(�Bi�t�\��8@5SN�-���Þ���6�6R������C�[ZVnn�&c��4<5UX7Q�#w�$�5Za^ZZѤ�2Z���^��}�3P�VH �d� ��ik��e�8v�{�GK<{�1ά��td3��(�/+�r�3�bo��)ssw@���e������ʙ�e�tB=�H@�~-�/@�J�o���n-v�RQE�A�~�v�����(��(�x�w߱�\��,m����&�}�*����H����oh&�|K�#tu��|�;��lL���\�zt�M6�מz<��:�)Q��1H#��N&p��ѣ��%V6���p���6����!�>U�(dXpw`��48:�G�P�9yV��Qi󰳓����%%5CbLíI<x1I��S�"�v&�$v��{_qH��/0�����(?��Mګ��^�$4f^�~�Y�Vm@G�0�D?�|b���R�k���tU�s�`{�r���a�3!��0��5�zm�jq�h�p����|��و�����4���1��)���Я�����ս�����u�ߦ56h��q펹��}:�V����Y�C���}�:=�V��
��;��ЍF[�㓶��;xٜ,�t�(�Jo��;�$��qs/��FXI�a����m{�P1�@U�١|y$Z��#
��v��+�5�>��ҧ�4��,�8�����ԍ�<!RmMzȅ6���f��`kl��]��>�t��5M�0�<���b？���v�[��-T�Y��5�|B��Nڍ�	�O��r��A��
n�O�����7�Oz��#`�S��O8]M���9���q <�묐��ń����fT�&�f�I�t&��d�{�lc���ߌoZ�G4��5��R�1�H�dp��
����x蕚�R�D�f���侏�㝗2����-%�O�Iӹ�d#,]e_�x#bJ�#0�L�39�z_}�):p׽%�h��0X��nT��]`�8s	J^��Wí�iΘx+0�MDd��ʝ�:����W��/V�aY6�����A�y����^�aUt�t>u��ɨ�h��l����i6�6}}�������;���//�~�e}��;��	�SPP�>�
	� C)}0.��o��x�D����rB��/E�+�7;_{���QUxE��U[/^�g�w�z�WcK}��Ź�v�L��{����洰c�:ʀ�S4�+�l����>�>^���t�7�D�]Xܒ2-�I	o$�P��F��r�V!�Ҧ���ȧ�j���)������0�r���d����v���=>G�k�Dr�r��?t���+�c�=p�%����D`ݐi�/�~��>���eŇ4�ζ=�A���'����g<Cع�ߏ4�lf}{��Q����6E��J%]������D�D��K>V�dD�����d1�]6�4��N3�h�h>���z�&��H�4ɿ��u�������7����7�X��.�������9��p�����⌴��%������`�O���?ϧ1s���k;�e��,���gߡ*���C��y7�b4�]WW�L�E��(Kh��[ \�?���R�)�rv�i�>���ل��	����Y űm�ww�����0H���!@pwgp��n��]B��5܂{͹�:�u�T=ӳ�Z���-�B�V�9��՟��Ȉ��/��7�`��w�O.�*z0�.��"ժ׍�Ѧ��v�ւ���xw�8;�$��Ӄ[���x�V�65��M�[�(�_�&�߃N�*=�.��E��yrs�~�L���R�uс�@N(��83�� �Q�b0��om�e�OL�Q֟A��ĥ Sڼ;0Y�w��񜦶�%2EA���\]1'w��(�<P1�����x{{�=�lTW��`1�?~$~>�l�ϑ��2JEgH�Z������Ǐ_f��(��o<��{�,Yb���Ƴs��⪈��/)��=t}I������Ɠ�X��s�Mb�y���"C�`UZ����&�W�ck'�h����lV�����q#�
h��l�pT7��53��Qo�����t(�'iW�=H?��HH}�,Jˌ[��Y5��eѴ�v����o�Ph�:DҼ%�%x+���aV҄��t�kU.&��
�ӣaV�B$NV$vmwvx�o�|I���VQQq�/�B̓y&X$�3�/�>/EKӾ�W^7tϺD1��=:�w��{ma�|d��vh[�'X�6�۸�����72f�vj�9(�(���T���A�n�$�������=o�f~�_$Y��9����UYj:�~�����jlĳY�NiG+pj��"t�ؖ*�o�.��x�@dy��9���N�yO}<a��\�������Y;���k�pM��;�����;���r�[�����z����(qȁ��#_����P��U(����n2S�A^_�'%-m�ec�6N�ƕ	��_���*L�p�M��H���:\H:j(������b�}�o;���z�?BM�DiV^�f ��8�O�@��6M�x)̛���KZS_�A��*�ǆP����6��
�sv����Z�F�F(�߆y�'v��E��H�|0< O�^�f���3y��ΫIA"N4\�bP跚����Jी��¶��t~��b�i$~��}�*r��=g�sMn�/���7��|g~�33��L|!��w;2�3�Ô�ЙHK���3qS�'+3���[�l���Ff:�/C�	YT�g�p��3�a�s�-�.�4	�+Kh_Y#rJ��=�xI��s�ȗ�T.O�ױ�`�O>%|K��N��;h�bz�܄%�r���e]��OhS�� �e��-�,�3�V�0��>�NI�I��ndM3y<�&|��wW$r�Hyh�F9�`�W\yԅa��)uϲ��)���l%;#c���'��v&xfX�J��VPͦ?��7��Ҝ~g�i<)e�j�՛�#h(�k����X���̫����Di�k��a����|>wl%���@<�]L�P��q�:�c�f�a�+߷�ѐ�\��&�57?�Tbd���t�t������'�۾���w��10��3�+��60PQ�U��SoB��O�,'�}�;�[����_�J���/�����X��,L�[��S�Kr��Y��'E�Q]a-�h�h�<Mb�U�/S]��ByS:��C��`L���_��h4�6�����t�@��0����9�Ǩ
��ǘ_���I)LA7ha#}���ב��{���r�%빏���с��\�p�J�ӆVˇoҬ-8��Ժ��#�&���ߵPZ��N�-�� 2AO�yP�lq4��&����DRM-i��.d�j0�Vfq(;,[1��o�NP�!�k�����I�i��K�n��9֛�~y<s����:�-hkx��x�}F����!'g���'�
r�+/� ΋�3^�Θ�gi�p��Dħv��裋R@j/>������ʸWߢ�n��Y�	� ��Oڟllr���@�J9B���EEw�r��̆&����;��G�n�T������K�m������11-Vj=\��C��,�Kٸ}]�!�bJ�I-`T�ŕ���-WRS�hB$f��Y)���f���9�}����T��S_F<=�ص��MA
 �%���>�'V�c5�{m�i�+���A����W�8���n?�G�fP�s(���}D����BW����8	���T���.+�FO��֌іDB[��Q���*t�#u(ˢv�A�KR�)�� �:����6��������$_57{y~RM�$DĤ$w_�v%����(aRA w,^�.���C��{g؛�q��8
u(�~5��N$ �v�U�A(��hA3vy�kA�)�|s�����*s�a�<�d����RrfD�R����>:&0*�����Yi�N25�t�ޝ�^�9�?�L��NiiD���1'����tə�	�C��������ɳtwC�j�D�����}l�F���Ϗ�����߃m�����X����W�Q]v�!r{J�~DV��bk>��D���l��/�wU�vzUm�5��qSɛ��	s6u�?L��,�������VE�I��<�<��.ڠ�$�}�z����P���C���U)���:_7�Ŭ�ء�� E\,��>����3�ĵfD+s�IS�(^�F�S_� �gec#����'��6��O	4���:��I1G�v���l�ƿ0�)�����F}��|�^X9M�k�?]��X�����@��KxxѮ��zp&aߖ|m�W����vA���iE��( kc{�t
h����ǻ��5��dHўK[�M�.v��ݮ�i�Ӵŉ��|�9֨�󛈫�)y�� 9P	A��������g������`�(���j��/Ա��Z�M'<����W�ߊ�����H5��$�%�?�c��G��^��$�|�~{�{���!1t��Ҷe3���蚅H�k�U�+zv=���Y�C�����v��%��D�%��  3
��uq+JJ�J �fbaIj��)���9Q]z�7��/�n���"�A9�?�y#���ö���[�oQ���}��,"񖫸���o�M�oq��
��9)�:��h���C��и� ������� /*G�bT#d,cjx(��ڷ�񤊊��A �CU�*�ª*�C�o���S|ߢ$������$�(@*�����~ܫ��$����?VWߺ��s|����z%7����Y�i-�c�GDל�ol�Z��(W�8R�=���#S;�I� �ܵZ�[bi�ӓI‘�y���0#�sg���Q4�!ИB�Ŝb4�]�������F,�*!r�d���	�[N[mׂ�ZZ�P�Wf�;8�����T_�uh���W-]|5�����`GVD5--Wd >OZ�#�z�a7���g��P#��Om4AI�>�<���cL���F��jV���+��7[n-�s�w�n�kid�b
� ���-��1:W&$�?^� Z�X��t��fu|���ϯ�w�i�ol�Z�B�8:;"u�4��H��z\�e��#d�m1֝a���?�>�|������ �9����г�p�*���濣�g��񌥹�mm�N���L0B>Ƣ���5c˒�d����t�' R-b�U0���p!b�Ε\_�4%�*����m�֔�)��;��
Hep5e�3'*�C�@���#��E⡳sr�9�\��?7DE�OX�W�/��P.��v�s���b�k'S�mr-�]R�ֆ�QΥW*.���~� ��P�b�e�;׎Y6O�̙�rˠ��0�'=N~�ש��%=�/����L�C@�|@���G7-��#���2��kŜ^�c �y[�xCƔv����ym�������n��W}  �jv�͋%ʱ��5xZ�g��.�k�Ɂ����N�?� �e:�U�Xi�R%� 	��q���h������B�� ;�E��Z�*i�^���QE`�o|Bn���qvQ�Ț$3��T�e����Mq)�����b�pӉq�V�m"�A��ʵ��gy��i�N�F$Mʰ�BIW��ڕd���"���s��$��^�^Mf,tH�inF��Ȇ����0UߓQ"Q�P��؉p�Ӕ��B�=n����B&����\��#�����0Z�O0�u����}q���*�;��X���GK�zW�����+��Gt�؞iX˦����͡�����Y)�n����� 5,	� 6,���)�
���:���2�3w`%��ױ���0���E���w{(䢹dGXE|/�"���?m��$�r����nκ�O�W���\�\�U;5.�����؉���z�PT
�}��f��d�T�Vt�ODN��	����G�v0T�?�SD������ (!J��3�EC�۩}u��܋pҴ�3|"�[�����QJpB�Pp�K�#�{�^jk|�z�n.o���Ͼ9Z,��iّ�K�w}�Iq7�ٴR�����*��6Ӫ�.�r�ѥ���7 ����{ű���0n�"�v�9E����S#3]w�BN�(��Ƌn���l�x���G������W7�P���v�3v��Ƨ��.�"T:��}z�)!�%{��ڡ� ��{[Ck>�D���JU�����W1JY�zvRy����w�b���	[�)^ ��s�<�&��ˏ 7�̎��Y4e����U45��H��E�T�����M���cp��>s��(E0j7}�=�#��f�|i mC��f�ƍ3��x��e��@j��Q�Z������묜��W���}43{������{o�i.8��|�ʄ���O�N���2�T��MH����cY��@��������
����,�Њ1�����"b�"����&
2r�̈́� I�@�$9����'a��ش!��������y�2rê���P�� �Ï3p�q�\���i��`�,^���ck}H6��=6�H��o��+ݍM��`BcS�t^��q�~���y���c�ˉ��(�+�j�q�vô�(烙�?~�$]1�Ac*��n 	|�3Ws;���fy�u}��D�l㶉yx��P{��ө�6\lx��1��6Q�p/+2.np�Y7)s

<<<##c `����%)r��BѤ��N���F�pT�B���E��h��s�����y�M%�� �G��+�;}�L/�~5`�><��=��Y��ِ�m�w��אp��ѵviE��<���'ojZO#��ݔ�Ѓ;�1��
�f���yУ��y"&��SacC����0I�q�n
~3RF�9xc�j���@�U���J��F,�mL/{:��^�%dZjۤ=���[6DVǺƾ������r �yc��Dx*��[�'n�H6#9��b���c���j�=�֚��.Σa��`�:CF�3t�L���m[zO��ի$,l�XXқ*i��-��k!���9QH��ݗ> �#��!�<m�38)qC�ѯW��]��o��F>�V
��6a��f(w2�R�m��2þESi㱅��Ϭ�gM�'b��][=O7H֜8R�R�8K������g����q���Í���OH�WE�H��]Q,��p'9DN@ ��#$'/+���X���2W�\�����V���ŧxvvG�8�D����s���
�������~Xq1�}66����p���:��#������0�=�ɶ]"�9�*[a��x��u�*ow�:;��/娱 ���f'� D�I��׆CG�ӷ�j񐉽�j�]�So����$j�/��Vr(80�����ҩӯ3�
U�,�X��(���g[7cxX��R..h�V����8��sJl�=k5|+��N��������R���`2�wð��
���L���-���w�ú')r��Ǡ��R7i�W�;u��<14������>�"w���D�ec�0Սi#�x9w�Ҁ�����D�v���1�CF�J���F�]��N�I�Î�`�}�H$[.�[�:D�ֻ�2�:^4��,�\l�F��������D���1��[�%g�;ZD_��=�YDEyl�`UPv.ŏ���<�/ �2n^|Sa}N_�e�eYv�D�<p��
4//`z�,�ﴟExi}�)��A��>OOO�غ�in� |���s�������A�>�-XFF�p�e|qQ�R��P��ɫ����jR�b���E�����fχ
	�9L�Y��!�1+�v��������!%S�M<���n0�L��Ur����]�����l��%*�	��p�t8m��k�XR�0,r|��+#fe�� 
$h�A8��Èjb�̫���N�5qH�<������ۤ��^�����@K~�28�\�pq�x���x�Q�}:���
1���y_~q�����| ������dc��цk'��It��c��_��L+�o�:�����
 �u����a���Z`�ւr}1;۱�������v<(k�+q���[���S�Ɲ�֢��5l���j���}���,�$�� G��T+���}����kҳ���������v$�i��c_��3�V���U�8j�,�Jh-�FH���ɳ�����f����^���Z�U�I�E��Ԕ���7:�Yp�)g��o�ռR�gJ�v5/�Q����I�v3&&��E�,@�T���s5�[�����x��'Q52�ڋF�t4�-��N?�)�9�q^����G�۽�p���������{Y�������+	i���2_ǵ� ��HV�gQ~?��0PL�宅X=�;ݥ��/����<\�/����sP�ddk�����W]�aV5��8RB��\�?�������_-�ЃP 弹�+��}�4@ʖ;�{Zr]9�
�$��O=�$t��],Y��x2�Dt�I�Ӵ@I�A�X���f9\AhV]�s6��H�X�kg���)�A�nrOX�e,��������,��
\υ��&���
�a{�b��v�*�06�D�a7갡�����T���U'�7Fj�6���m�{��Y{�e�����..���X�zi�p{ef�cT���p�!���U
f���Ūkwb�ֶ�d��E 3���ԲY���.�ͅ��?���C�����ył)��������~�<��r='�u�K�N���˛{�-u!�w��
^l��M�ZdB��1ϙ�i��o���	�v��/Q��F�H��|Dw��Z�Q4[5�p��ugp�+(k�#��v����������M�m����:����L�~x�ej�S��HE}���Y�e)�b���W��}�C鞩j�����`��M.�::�yR��C��U���eB���f�^��xSN�To�?k� �?wx��#=�j(��Ű��j��i��<D��T�<���s^뻹���w��c�Ou{CB?+:�r�&�]�S	�O��yX��g*ޫ�IǤQjr'�7	:��Q���JaWUU	�d`o�-[��oH��淞,ftS�[}e�Mz.tΧ�M�`��}�"߽/�l��>!!���Ĝ��[�4��&&���a?~��166Nt��i��ޮ	{q���B�.:����G�L�J��y�)�!'�y�wEkE�zC�|4�c��fYE���ě�	�&q� `�D���%��'vM��G���e_�����)N��%Xzk_���������n�"�S��*PC��=_�����# u3(���?��-���_?£��r=�#� �����t0"8����S�o0����	Xp����\����u�ݺ�.�oR�,���vM���ɔl�����>/���H�;�2����r�zm�<�nY�L,J;���a�]niv�=0��}JG��ڿ�۹�oXQ�K������)g�el<�o3me2�/&�#^ۺ%�����ku�6�A����@��sE)Gbɯ�{jk0�`���Kh�D��)�I������`�N�r0��(((ʪ�AM67|�XpѤ�v��8�׺��,����*TLo~�����,e�ò���D�F�/V�L�����$ߺ6A�hb���츉T{��y��
U����n�(X�����v&|�7CR���������R�qa���vi���#D���m�L����I�:R1�#7�6a�a�b$?4��3�(F-{�hK|�̵Qr�� ����g�^���_+N�44�l�Y���]�	�y�	���P��P��fOn�F7x4����h����!����J�RL��D鐶`Ӥ����l+�����P,�W��ʗ�k��)��:�S�c6n��*������!e���,��0T�q���<ue_zD�u�D�D����ww��-̏Xa�9	r��ݳ4E��������ĉf8.e6Ӑo���M��g9��יc�4�J��R��U�\����������ht�4E p���vLDkG�/B����*x����T�k�226�R��f_��"$�\�����k4hi���C�[�Yp2P,��=c����n�����ޘQ�ѕ�\���S;�
�N�E�W`��L��,6 zaz:j���u ��6������s�Bm���FE3l�~�!pa42�kM�����&���jph�ޖ������2��?�(^d!���tV���fl������o��B�XK�74��ss��m#��9Q%�
�����-�&Ƒb���x�ߴ�2��I����ڌ
N�H1�ȩ�b9�~����\5��eO�]�75��U��r�
��>�G3��s�[���z+����=TR���acji��l�e�:E�����?j$��Rq+�.��L�������:L�v�8Kw���b�"������t@�өfU/�ׯJjG�)�fjY	Q�Spr$:�U�)�{_\�x ?O7�u��=��;S{��V����x�"` *�l�r�����F}Gt�nB�2:�4��F2��؍uU�n���"��?7����͎.�ud������3.�!�-:E���Aq���`�����"S���0'�0Z����?/6(Ϥ|YYX�M䄞]�$|�����5w�� ���a9�/yJ��S���QaU��$��'6�<��-He���H�vh�ԯE�|�CY���9ĩ.��
~f�E������#v����إE�?�f��k��k����p�#vM�ƿ@�OiA�G�cz��ވ�X�x�朦���������:͹�^YA]#���SM/l�����n�[���Q�����.���(�r�[+db�-��
l ��n��O�{���d=&f�N��G�c�@�F/Z���M��*�'��"�O��������m�79����ӂ��7�U��߲�4��ŠB�ck�
U!��
EbT�0>z�p7�ǨݛtX������Z��"�0bi�����>��~� 2���28T�[�N�"��W$"k�cH�M ����:�3���Y�z��BR�!�4���]:l�#hj*�U��A���o3^��#Y��?Ԃ|a����Q۪y��K��J$��wg�:����=�s���L��M�!V bi��(ee��42�G&��\� U�MTS�-C�fn�WW,[���y�Q�\����6~]Cb1b�,�\�6>r����"�y�P����9B1�A�$���'�=�
:�v`���*�l<����4���ʨ��g���[��/�9/�C��#!�����K���ޠ9$�T��@�3�"P��T��p�/|�6�?��6�E\{	x�����=��?��q�5P.Vެ�_�t"~h��g����V��jX��U�DW�C�8�V.0S��$yT,Y��l:�r����0N1���o̐[O���Ň�J*�J�`��;K7�7z���^�����^�ҕU�`P�A��P�5x�L���p�������*����i\o�}���`)턁����z޿ɣ)�aZ�
������
�Ï܍/k�Ӱg���������U�]\�S��r�s��^��g�0�=�%�ǵ!�,9��3�P�lȱ��^�%>N%x-x�������>��LE�����\�����=R����]�W�[���U��eX�<��P��iG� i����3F3������u �U�YQ.f��Ĵ��e���B��[��mj�#�ED'��*�I����گ랪=��EO~��<��6`k�5�I���01�v5�h���§�U���h��P��m!XrTy��o����wEIu�M���҇���D��S�p��rS�N�;"�p�MDG�NiMi�)�Fn��}�w)S�D�I��'���wo1RlZ9p]~Ȉf+���_�3u�S0J�#���7�^�����$��D��>b�����h5��ņmll��C�x�~�w�a�< &����}{�ܱ|:�j�v�B��f�
����/�\������vs���\y����R�� �Y[�/� �E+Y���97_���P����;�e�U_L�v%T��b�5��#�sJX&�mzw������f(�x����1N�Gf�c�-CCE�߻]b��M[�߮|�!�+z3�����ISa�9����$�㽥�U�ޔ}}�>��;O��1��CCB�}���0%+�|h�E��+9PY��Z;1r��v�Q (�=��'="@�Wc�������[�"#���od��田2���M��p++(��WW�
��-��[ol(=��G�d
����p���R�Hs�����^~��]�r%Qn���/o�a�.��)f�|7�Q����؋�/VeFr�F�S�m�29�����s��]C�I�<�q�����{�p(�^i v�飸Y�J�N8�����f am�.Qi'n�˒B����e���P��p�H��G�7�Y_��n�}�<���![��·���lQtÕח�'��0����e�@ֽ���j���p����b��p����Y׭Q�mVW�j���If1�R�n"����s��E[��I�~��squ5~�{m �j�/�.b��w9m�v��U��ք)gݯ���1{���0�h@�a7t�֎��GX���>˚ʖ�SƄ�ؾ�5�oǻ��
Bs���P�̊sp��%�Ut��v��|��t�̉��2���z�&�bG|�$���x&����6wd�n�f\�Wf*��ʃ}ȼ���n�	{�+$��sp�i������1*�����K���jv������q��q�a�L�j�ޤj�~��}����|��h�<1{� *��(qC����<1�ܔ �tzF*����I� ���4 �Z��Ts6n�N��!s�JW��<��X��g�ee�x�S3B0ǻ%+�%�yQ�q�ȁ���b�R_�����l�~ �\hQ�RMj^j�6�i^�Ÿ��[��.��"�o�ނ~%3�{یtaGg�ka�L�Д���A�G�j� `G�������{�Z�B��̆�c;S�C⁑���u�do"�Id����q{ S��{�{�]��p�XDP�D~�$�p�~�?�	�<-�\�Sa�H��o�/�s_�h߄�u@dI,mH/��G.�(&u�R��E�o�b����l���%�+��4U����@���Y��+�)��N������\H�o��U멲3�Sd�d�L�;yQzA��쌣$'��/a�����u�B�"L��U�H�e���Sf�y��4�X��͒�_���c;$�7�;���P��rțɘ�1�t���Р�0|�I�l�;�w��=��KAZ=��W���Ӗ*�m&Rq���͖�kJ���%��p��V��U=6�={����ޗ�~<Ɛ�	��?:��Ŧ�4�&HE���_-�|�Ӓ����K��#n�S�^�!��n�]��^=�w�2��v�̗8�ʃ.�0��S�J��)�����uܖ����Ohc����������r�ӃY��CD֙�G��7GHo7	_*�a��i��3�N>SQFL�$�S���ҫ>�x����4��wwB��TO��	p��Ѷ���ZA�l�P���"B�ѩ3�W����׫'vfq)m�{�w�n���h��mqI��R�y7c�l�p4q0 7;���~�6��*������Kc��}�Ĝa����O#�l��؜��1�Lx��B|��ƪϚʫ	X�ڍ|�9������-�Q6��rܬ�,7���Ȉ��F2/�?�*�r{J��q%�	3�o��r���*E"�5E*X\Lj/�A�uЈ�b��Ja�Q���|�V	����J��b�Dp�!^�4B�t�����I��q^煹a�N�ac�l���Kh�����r��	S�:�1��[�b=�e��K�Z��W%_���;rh��_������'Zi��X̀��,s��߷ �nΑ��~��#/%�V0���U��E�<XED�H",��$�b;�f�D��CXD;������5�/�!l�Wr�&(��� uè5�i7p�K^������r����g�)�[&�w�������,����D_�K�� ���s&�G�J}s���̎�I��
ͯ� ާ���=�rą4c�U�)������Zl�䩿^������?z}�q�0�O]�k�%E��!��J3�4�����S�l�������c(2����~=����{�f���n'N���b������鶰��>i�f��|`�����d�:�DXX���e(۸�v��R6H�nY��;�����9����=o�B�2���o���x�|�;�i�$F��I���!%&�j��Q���g��g�~�s6���5����@%7�v�	�Qӄ~�Z���|��X��%�O=Dɕ���Nb\�v�_3J~�@�ʥ̜�(��.*���x��<nk���j�܊ܑ������N��~BB���jg8�ݸ�t�=>l�qOKS�b��)[ZZ��9z"��OOK	z�Oόͺ#���T�g�hnn^�w-�	�����ԛ�""/�����;���]�C��-����Q�٠���Z5�k���~��2�r ���w����Ɖ��K�0TV�V.h�����P�F4��bOf���g�c��<�����0��c�P�nb��F_<�ӌ�tן��[���U��)^�h/��	�q�.X�B���wv�%nU���~ �$rH�KN�:[�y���[�S�W�9��D?������:%���}dKL�{��"		�e����"�=q�c���PW�?��u���6��
�.c'X��c�v}�	v^����_�.p�D��Ll'��<�
�bLq����xʴ<1�=.H��.<4�kp�Y��:��fq0��qc2 ��q�9��
I�1�"��F��'�����-�׿L幰wr�i�����X�PȄ����u�JYAô�M]F�m�O�T�θL&o'��p�а���;׫��
�b#����m^,�b�#ڈ��	�b��o?���?�x�a��<�Z�%fmF�g^jb�ɼgQL�N�sad��Z�ի[Lcw���M{l���n-��O!�q��o�F2�'=�Vi%_�N�`�X6��x�d �W�0Xs'��b���"���W����$�@N�
���0��K2I\�x��>{9��ߊq��o�AD��F��_T ��X��<|�}'@7�ث���;������/4��
方�.˩�3o����Aj�0��z2��y�-8yl7[�IHI����ً���6�1�x2��- �Mp���Ml���E�b�u���a�̘277w߁��g0kJUU��Eʪ?��5�j�� w� V����ۏ��f�|��j��$ s��g��l��ƽ��QJs���IDF2��k�Q��\h���[եrOm�c3Ė�ֱ�=�xIZ�\6�n2�I�tɉq}'
ɇ��v�| �?�����/���9"o�\pd��o��~Ib2���j��!���>���l��ʮ�����X{yM�)�(~^�a��_�+���K��3p�͚�X]Q��6���t
�X�a�_w��r��AY\�;4oG�a��%�)�%��G�(Ԫ0����q.��LX6������6sn��y"Oks�%�n�DݯR�y~�/&����r����ru)���Ě�}�F=�$�yƐ�h2���:)ҥ�V�v��5N��b�[��s!}ű�q̺������c-�x��2^��&¯Y��Y���6=��[�Ys*�E�N��}@�KT=��̰ݢ�yo�g�&C�_�<�|���jo�kq�����mS����̯K׮� 
>�������!���"�\�m�����[�a�ා�.!f�?�޷��x�߬�?�zT*ŝ�����\�o�r�\�b�9j�����;�v<�Է�1`��/��O#*�V��g�^�SA�'͠��+"�EO���q�į���0E�9��x$�h�%��EP����E*"�8�G1�@��	�7�^g��=�f�?�A��(4�v4��S�¸���]����m�2	�I�?�)�c�U%���|/�s��&�H�#S�-��m����;��4p$]l���x����;���:�6cdo��g�E�����۴=��p�}��:t��>;��c9���"�ץVevȶe�����9I絛���=R�;~��6�,�P N	(L��M" �-�S"�a�4GD�@9��H�ӧ!�.�v�%�yH��bć�0�a�a" �ޒE����
j�U�bUψQ#�(נ����`x��H�ĥkkuZ0}��� ��9���0f���(�7/]A�����g��׋��T�-�_����<���g�y';������}�~C7r��4��"�^�����UB�.�賎/����G�X�؁��-Sy�F�
9�R*�O��b��,�n�Rt��*�2��H.�jC��d��8�c����] ��y��dyn����4�����n�g���ͨH%QZ�ʰ�1p��<��۽�$�qƓ����׍�7�ݏ����3`�IޤID\F���JKٍ��%6�'p�dV�����5��dα�GS=��&ە�W�� n��#}�	Y�v��M����8p�{!�O�FV�3C�}߅�R �e�r��f�!N�؞���5;���=�k, �]����y}u;�̗;_���j��"  ��<�y�p����#�
��ivbԆ� ��C^hX�X��{ 9J���=��&H�����\"Z�-Ŋ��M��V66��y
u�e��ع���U?����S:���d����o�:������2��O�Z���`�о �[�z�i0lt�������,#��uS_vv6[愕�}��I�֎������8����	�RR\)l@ؾ(X��I�� �%@4���t�.�.mzXR�$1Py�_��欱IH"�P	0b����C���`�7���ts�����nD��c�������-�ſ�>	�T)[��r�7��m��vmo�5��nf����}AP��2���$�T���������%����1��_w��m�ѓ���ω�vࡖ��=:���M�s[���l���[���(J!��g����,Ǻ���g�2�VW"�hғ�+��a�ǖ�b�E>�K�Pǯ���e�/7+f�վme�b(����Ż��ĭ{2ƿ��au��;�`<+��-�^�_,[A��+�`�܉����WL��U����$s
U�QDrK���ㅓ���d����Ã˺��-g���kX�_NR85)�V�@6�$��miD(�F������;� Eij�~�J<d������4J�/�./
������wS�l�|ȩ��!KS�꿄9˞a�θ���s�����>���44��7<Ժ���i�j�8G���(��
d�߻���8]Ջ���~�J����Ԥ�xi6���;:>>��A(0=�(w�M�?[I]K��������$�u���%C�R�Ԉ#���9-�scccHD����ۂ�,|��o�d��%�k)~�������4���u�����w���[[[�u#��;�3����x����~��H(�p`�B�F̜?��.y���~�d_.iu&��lt�TL*9�7Z�|oan�8'�^�A�b:7;	f`!����K�`��/'��Q�^aJ��׭����h�kCy��Y�h�a7O��Ε��7eI�'���o�Y$��3��V�P�+7�}2�����#��?$�]I�ɑX���%���nT>\�k_�#�۱)((��CCF�:]kCO�/2�=�aj�"�.�J�lB �u1׵�B��fL�v���t�^<��LR�s�0z���TF�!_� ���E��vm�
�	}(����üӣU�Rc1Xw6��j�{�e��������ؼ���[{�e����;��볦���A_S�*�����&�m���Ӷ����-���h�0%...�o{�NV ������tں��z^��l�O���g��E��?>>~Yy���3�����_N}}G��?fgC./��P~� VJ�t���xsH\�-&&&wg�P@|ܝ��D]-��Ofc=��*��(f�y�u�Z�ǡ����ˌE��{�\���e3<�<� )��>d�oR����u�E�Yj�,d^Ɵ�^|�W��/�g�W��F��roZ�k�&ZVTv_��Mw�DS@�("j�Y�_�4����qu�25i���]�i�-.�a����R�t%�T����t���oN�7�#ҁ`N�ܕ�����:x��6�y<
q��NE]�h��z{܍�'9�c֝d�JuQ�ˋӛ���X�l��`��4P�n��~��i5W}��`=�@�s��.�K��𔭚&���h�KB®�C9	-ϓ��)gmՕ�]0zT���p�v�/l{�D.�O�%�|g�Kh?%�x�ke��(��LX�=�%��5�X���|N2Xu������K"c�6�������+��h�u��u�@� `����:��@���݃�[pww�5����sN�bA��f�k��IUM�Ǫ��J�8օ۳��G�pسی��P��F����ڕ��{�]��8�@�JX����1��8�g��n^�2=�h�O.�g��P����>F>�'C4���z���F�|��*]:V�f|r2 �.���H��RqVU�L444l��0 1==
.b�����i��54��A�G�$�ҁ�<����祜(������bfzz��≭�&(yh�nH"'N�:��KJ3���T�L�N����cJG^���ux�u�p�y�p�
�C�6W����&nŌ�KM��K���kY��	�j����E�
�����:U��"�1j�Y`��UpPj}C���h��hx���[+1���@��QԞ���!�*���JI��նk��p�,���ܓ�y��J6�B�����.W�d��<�jiDf�+␺����2���7�����)y��.��l�Y�a�KM?�`�����B��ۖ,u)�-�"d��|�UZ$�ۥ���E�l+K�&<QA�]�Vvԩ��.N��&�Z�Gs����\�\ŷ�V���(]�I�đ��R��?i�p9��{����|��H�����x�ĀcG<�`�?[��\\�����E2��}]�\12Ft0�����`U��2�E7��	Z�1s��4��#�a �g]!k��HzZ�b������I�i��,�oҩ�x����	C��!����:-����M��@@'9 s�*:��}��(𨗭�g��w{��Nf���E��ˠ2�������Nh��������T���w&��#vqvU���t��C�u
�#���d���':g��xKY΃s���>�Wb��A&�<c12��u���7O��Ѻk-�yĞW#������bQW�/��=��I����{u��MW����2)dr��}Bxw�b�S�W���H����G�n8�P���멘���s��|�%�5N�2��n�2���e�~���J�a�p7�ai�|��D���iV3�ي�y;qq��:%�mM�2B�-��v���i_����{������T@�D�/������6�Ј���o��nm���I$x8�EmJ�c��0@��������_�H��3�q|~>T����������|D��ɝ=L"�cg8ž��gvv��5�2���Q�MC���FH,6L�1kw�n��<(YFsL�����Ȃ��0I�r��BA/By�kӛ��Y���#��Z��9t5*��s��ӧa��G驯:c���B�̲���ŵ2G�GE�9�cOu�[�d��uz��9b�ap&�p�05#��^:O'>>[���|$aq�o+��X}�O��P��h�Q��$��s�Z����v��o��g�"/ ���U�\��K�5*i��o��m.2��4e�v��;[���{a&9��`v��~��z�r�X����߾A�,�>�VO�[k�fR;a9�[�m���dA�继��]��>�J<���ݜ�N��xn�ZaI�:C���(K���S*W��s5��L	,��wDD���')�7�u;P(.I�#	�!�?C��������k��;���Ml���`�ӓw���[�8����{�)��V�{����ꥸ���������=�()���|������1<� �lmYI1�G#���8K�񕕨��욚xTŐsy�dޏ�� Zgi�P1k��E��u$��4P�n1����-x6�Ե��~7`k�t��_t�C2w����*�d�X�q�����y��у��Ϭ֜iA���[��}*E�g����m�������~���o�NL���FO��JR��@R�����$nsȣ0Kk�\����y���Q���~@������w��b��h1|��w�{�?wΉq�0/3��zI��p�)Kt�aۙG#���˾��@���2�+������tQ��+:6��P���P2�֧�:S�x���Z���[�U:�W����#_</� �*�8K�-�]m�ڍ��d�?γ�M'
�:"+��OI3U�돉d����J�]���EM��^Sq��6M��G]i3){7\;>����܊���$2\qX|3si�c�8�r����*�й ,�����!���_ �@�@ g��-��U������W�HîA�?�ҿ�ېh��6{W�H��o[-//���V���d�� b(؁�Ȼ���o6��pB��E|�s���[�3lEE��"qv"�g+���N�(�o%<���b�((���;V�࠘<�*ǁO�S�/ZzS�X��y)
�|[-� �T�A�x��YW���⏘-�����5�ɑs����DKi�c��}	E��}�ܐ�s2���͞���hoӓ>J0��˵�H�[���.u��K��x��li'ixۉ�֩��#�t4q��Ob�U�������������vՀ}킷�/�F�U�϶&WL�����q���5"�~����)�ƭ�tݣ�o���}�A%���=�Q��h������foo�q���{䊪���DH���JT�ʗ����I�\]7��(�O�hW���A�R,��[Z���:����d�կ�֫/�\hȅ�˗q񪆆���=n�X)�);>B%�(��ndkkl�Րi���U1��ora��M����8���bE˜'�X��`#,����_1����D����ۂ}
�����W���L�Nf�!a�12�`-F���w�������
{�f*"�+V�2�'�P���sr_�#i͎h?�-^����/l����\ePd�5�H�KF& �ĕ;�c�P�$SfD	�����~*���zc^����;1����.7d�������nޒ2
wP2oG]���(K����N����\�x�, ;��H�^�r�J�;���_tG����g�d�Da;m�^��n���8�8]`�ױ���qm�R9��K��k��l���4��]�g|��y��"|��$g=7V��o"b����
ئpY��֍��1 I�������A�`�R�0�y��~n6Ļ�����˵W�jٍ���	�f	~�E`�A�1��XzP�TA�����Goƴ�p�'b3ҋ�4σ ��)tK��g��&[�6�cq¶�鸌�B.o{��u�u䇿G0'�e�/%]i�Z�D�yR`Փ�@$���h��~�ŋ[#u��[��j���I����2b�`�*��lW����4�.o{�!���}��#��ku\�6Ghx�_�r�>Q��m�.�}�uɲĂ�522�s��swwYe�AB
�f�R�C�T|�#PcS�K~�3��e�ѐ<x��/{f' '�`�+�q9��W�CP�3�������Vʴ�� `�B�g�s[t���W�p2�7�1�?�qҼ^){P5��	\'�'�HաhZr�M6���qH�������7�|?$�v��	�y�C�,�d�j6�R9�'�'�t��}���f���i���553c�M�����̘�Xf��!�����^� ҄*�4[�RNb��c���».��+��E��v���w3%d�%���N�R��nC��o�ez�
���Zچ���+�m��^�>=���e�%�-��M�~���9b�M�������#��OuB|�7� ri�����%z�b�B`g[������U����L��S�7�mr���'|Y�{z����-��繸�����]� �:���f��Cʟu�S������1+���ewN�x��%�(V��E�	^˃�ԕ,CTS�jY�y�s?°�5%�7��'�x��T���@5$�q��xS��O��I�Z�6��Ӹ�B��7�TQ�B�֯�����+)3�}ll�d0@�`*��}�k���Ȭ�I�mG+��ui�.�M���+އe���YLCX�k�J���ӯ���?`N�3��R������Q��q��ed-�ͧ���DV�}��s{2w9+�̽�C1W��V8��.��=`i��N&O��(>!������-P�ї�l۱~�X`�B�N�����ȋ�R1��P��?�pQ'��Z�t5k�,6,:Fa�I{��}+%�w�^�k�� ; x�/P���w� }��8p�P�'�)����u6�f���N�s���XY�e�k%e�(�
�5�,�P e����@�~���Ⱦ*6�D"E/V�u�T��}���̝aMo(/5���������ui�Hؑ���C���w���Ά��0�rD�t׻R�sU�<������?q�;�_^���u++g�(�.j�z�z�&��%י%Y<���1�g�.���a��b	p���vy�"{^�z�^ۍ�,55��X��OoQ��(���|�v@��)9:* ^C�h��^v/OP&X���G'M4Ws���m{����@9j>���� ׃��/~'�(��>�N�x������,~G~db/?�Q\��;�q���Xs{�O��}�z���Y��C&П�?�����+���z-���\Ĳћ����v*��������E����>��k�����.�xc�G�a������j������\>�t�mPϥ��<j�r��2��|b�}R����U�G
���~�0sݡ!Zz���"��;l*�|�]*�M�>S�9 *
C��Q�d_\���k�65�@�S S�K[�b5|(�����Z�xMq2E4p��kt�m��i�T���'gA �;T���t67׌��a!f.�SLp�O�Rdχ��#��8�����X�	x�*�lh�����|X*��px7R�*6%��(�b�μɟ��v�9�
�D,+<���5��cEx�2�!4�gr��,B�
��J��_~�7�>$��I�����RQ1hP�W�>F
��K�c�E&^�4a�^5N3��x����6=E"��1���ˬ�iA�j���",�VĈ���U���{r�V
{���ݸ*�5�,��ڦ���$��mv{ϘU�J!e��D�e>�?Խ}}�(��7��:A�8�;š�m;lq �?G��X�?G�.rԸ�߸�gg��{!�a!=�5�]TPAdd��Łæ:,}���+n�d��׆;�Z2���@�Js����Cи	���n���Ӓ!Όs��@�J�� pi�N;Oya�����kN�a*��4�2.7
k���Pz�x1�i��@�����	�#���t�:\l�u�:�&ȕ!�59�{�1��C�8Δ���i��ȮY�Q�^s6�`P�K�E�׊+o��U����`�|	F|��F����������Y�a���]f6����mW麎����i	��ǕH]�677횖����&tK��~*uL�+��g6�L3�����2��DJ�k��O��6�X!p̤�A2���3ZX���_ܝ-X�g����X�K��������w}��s�rx�͍����H�����֒-B��R`��#EƦ�U�b5hÂY�D="!o����ao��P���8��]T
��R���ED{R��s�>��_c�`�Ɇ-�����c�d0E�#q��7��U��'
��+K�]J�zyY�~��<��iSi�5�*��r���y��J�A���%C�Nw�gBN���O�=e����]e��H�1!����/� ��06�)����(���gK���"&�]��G�$[h:OW�q����$尙Oͼ��@�r�5��u�]p6�l7%^A�%Ml��^>�
s��|��&�@��Yˣ���U�F�
�h�v��5�c-�'d�l�����C�8Ê�A���A����s��O�(V�Z��<Rf�-�}(ؿcFN�ޝ��34����"⨠�����I��Ec��!�=2/�������fpς����>3'�7@�-��l�d��AI6�O`�>�3ܐ�b���\;�f15�z�y:�R��o���v����g��y�܈�P�Py��#x5�x�N�Oy��B ��y8����޳�㎯�2�x/��+�4Tϑk��/l�����q���������'�D%��A��426���,Ysd���YVd����Ej.�T"�0l�:
H2f9U�;�x&�L�mZ-�ӻZ�~�
�M,@��@��tYf&%<��1�_fo5d'ό*�c��!5��@�9 �\��5S�ҁsژ�P3�P����tN�X:}OM����W�?�y�@��=��Z|�PoX)ꐽ6J�[��Ԛ�uN�pH/7 �s�-�0*e
�����i���E�Z 2���V�����0Qy�d�V/�
��Wq�Ҵ�=�p�
� j8�B�^�Q�T���}�r���es�i��e��[��`-�>@�y}Wf�ҀZ�Y�v*`�ϞtK<#M��̙(�"bo�	D�3�2�;I�H���/å��!oݜ^f:������9^�r�����u}��dV�E�S�̾d.G���w�R�Y�a�0��O�t��Z;l*�3
K"�|>�<i�҅8M|��Ϯd��S+єi�X�W�%`���7��J�D��}�ԧ���sBh����âʓ"�G� cΕ,�	8���Ǳë�}S���._l�;��������=,���54hu6p���3.r�$�� Կ��b�� D{���0!a��3�������p2_@���]���U-ь';~�:��\r(��o���G00�5E�hj�?����j�m<��L���H������D�՘j{�؞�®�;��o�e��:C���I��p���1�t�t��CX�B����Yz�!�n4m��������ܘ�8uL�/kH�u�ʐ����᫺w$���>A`uU�9yM�� �-�.���1��ܯo6��F2���5�p�̝�\��0�J/�������<b2('��{N��B�u�A�������R?��:�w]�Z����箤���ѭ�At�ߌnN�������R��BB
`�f� 8�. ��>�0�P�	 ����Tl\��W}�,.�S*E.[`��Q��TcN�� ����l��ar�^3;�����k���Z�6B(��f~x?M1({C5w�C�0Hoj$Wy ���F=܋󙩐xE�
"�jK����>��Q����¤zx�Ð�O=Vrq��们���WH�����ԑ�d���-���5
�T�HvSb�g�&�lo���V���Rw�K���TAe�Mo�	ׂ]_�H�z&n �vb��2���Ԩt�e�����2�O�Jō�B��,�qx���XZ���_�q�#"#)�dw���E��S����N�9�i�"��y���_t���9Oz�5{���JhY���ҹ8�=�F�����6��5� ��5��^�$���W���]�F�_��8܏��Z�-����f��2��@�I7vq+-C$��+��� �n�4��jP����]|�^̶��f ��}=D��b�)cnO�0w_|?>�C��}˸�w�/��r��^��$��ssC>:D���W�)��N��I����+Es;��L:h��P3~>'`fg��A��y�d��t{�\|v~��NF�F�&VJ1[=S����z�a��������V��,
E_���5Ӽ��o�^��U���?O��Hd���G<�!���گ��q����j(��y��v��Z��	 WY�Iҹl\\_͹�M��ֶ�z����;p���S�P��,{X���ZZ�i.v��4'�G6#�Y��5��̇���?�
��4.H�������ܑ���{(�o�J])�Z	�a����pk:F=ۭ"wO&5s� m��
����:�q�{_�zT�|�s!�7��oOx���D"�\.�.�T�·>��|�����LH�����g�8�qL��0�a��J!SRR%���?L����ե�,�[��mg�����R,P�6KkZhɉo���ȍOxe%;|@�f�*�m�M� ��� �=�$kc��M�b%�"ڗ�B��f�7�s�y��+p�.I/�'������Y0#��yC!�t�/BH8z��9կ� ��c�v�dS�3�]�ׄ����2���z��ώ��x�H��{<��݌�Fɗvsfx �Ix�~oȘr�N}��e��S�n�F�����E��6g2�T"~RghȐ�0�ߏ��u��¾����m��t���H�s��52�Xj�|hϰ갦�H��Dg9�{�]�e%��]^d�{G��q�4]� �N��A�9n������<�����s}�*od��<QKL����Rf9�R�з�����&�15�J��� �H8�K͠��K�&�������=j܏D�,䒏hD��g�n{&��$-,-���������L���7�N��[��nV	$�`Ҍ����{E�G�:e�ʡ�.��F�ﲀh9=��1�W����R��w�^tl�om7�I��ٳ�l9L��0���*i�X�l|u�y%�}�V]�\adu��z�ꚪ�|ܻ�	 �T1�5�����k���C�EK�:����ʸ�����b8
}uV���n������qeb>��%�`d�����P��A��~ȑJ�Gh��tƓF�'RhIV�q��t+���8����1|*��g/���{z���v�+,�:�01�D.����lt{w؇x[���wc��X��6ܗB���
���y�kS'��-�ų�f�~��a��` �ϋ$����?�-�w�v:��-��/iTRO�'�7NAc6xMU����s�n�/�B��cx_�	��U�3d����tP$O��(w�h��;`��]�~��fWC���@Q��s���j�_.������ mh��~��X�Cǎ�`^y~ܭ��H��J��Y�yĵ�O�{\
Z�:����uk������a�6=}c�7g��sB ���F���+��E��ն�Å+-������M�$Uw�ʏ՟�u=�� �xE~\۰��Y�;����{�;[\��ϓr�̊�=��;��B����׼q=]j���j�8g$�f�x�':��0�0_-�δ���� ���L|�`Qٕ3��<&.����%�-���=��^�uǞT���ؗ����s�*e"��Z��

��&��7�#���Gw5�f�ϩ�s�؄B�z�I��caz��n�yۼ�鸱��{�)i�������*����F*�d�̜B���RS?_x�b����7���QI��J���9I\�O����+1� :Z����ꂁ��W�g�$J��;��@��!��ն�`4$�P�-&u�(���P0\�4@aI���#is�^GP!**�� �t�"X� n�����bÎ</��uāb����jh�\n\�4�F�B�)8s�=
���������RK ��X��}ތA���I�u΃���h���z9>î���-*�s�M��oi2�=��X>M=O-_q~��E)�vk5~@E�j�zԅJ{�P�W�=m�u�2��)S�&��\���^" ;"�
�a��Y�?9Z���G�b�z��$S �����?� ���d�^b !Cr�(�Mps���/����h�e��f��2^:��R!r�Ńw�"��gYK�6��ņK+\�Vc+�"���)��e�Ї�ܔ�VX�+�;wD6e� ���tX�~���ʬaX� �{\����MA��~�(~cuu~*w���[ �ݔJ�l�����_#u�LHD�D���*Y�n�����)Mq O��=��Cz�蔂QZF�1e�A2���eV�f�3�Z�*��3�3Ox��gʝ��|�Kb��RF��p�*�ښ.�����T^�UN~��D"�2f^���j@�[�>{(KС��#]>��l��j������%)$�|��Z+ ���z��c'?#�C.p���b>��:��2�s��t�����t�/�~bEM��c�@/4Ny�(��K��J�	�[�1Ym^����@6
f�r��Q��W8sF<)U2һy�l������ Y���B���T�9��sbՇ�p�̮�>/K�=�ׇɛ�2o▓�/)�e���v��`j�|Ͷ&�Zđ�v}��A�D���x#
ⲰҞ��®3�*L�����0���	�Ȳ/�����3�V��V��x�[���\��>�0>?q�'AX� S��g�������kE(�*Ն�F��QѪj]}�R8YY��7�2���%�t��np�7�Wafx�F�~pY�����x!uH�[���J��C�f`�E�9T�ۗgCl	d�lf�����#���c###,�9�_=���&�+�4�kh�~{���P>8�ݿ��jjr9�*���GW <[EF�C��
!L��/5�J�����x�N4��gz�a՝�d��J]n�
dbJ�.�}���:;9Y�z��hu���/�*$$%c~�LGQJ�����\Cʶ��ge�M  �!MPJ�N�*�nY����u�nr��<�A�s�g�p��m�P<�e�:�:����K1���Pg��.Ha�: ~D]��lr�R�9T��I.���f���61���P�beV��x����7YP]�nʐ�c��f$'!���.�ҹkv|css|ǚI�e�&��e�좰b���?h�]|\\Q��5�Q˭%Dzm�4=��5y'��B竬���#"&++�ۈg�¢���ʶ��_#D�U\Z�md��~H\b�y�T>�%Q�U��W�E�/�+B�~����k��r�LId�c[��DL3RE�_��f�#Q�0 ,Q����w~�f| ���k.W�U]���fS���9@#�>ѝ�m�_���}���'�̈��d.K������Tݼ�֜F|`��S2Uϧw��$�����,d�n󺕗25�j��,�9��mĺ9Rl^���~��*d�h�2�%'��=�V�	֘�}ƃ_�����p��(��O��pQF�V�@����z�WMj( 6�+��"����8�$�9S�Z��+�P&̹P-�XM#�� )��4S`Eg��K�L�K�w��t�&B�z��� (A�ꩤ�*5g�QV�~R�![�����˿w�%���l>�;�X��8њF�	���kV�H�710�.\�KQ�m��-Gj�s~���|�Rt�dB���?pqt�G^�����4����߃��z-V�6��Ay�Ӟ7�T����o��P�|��������}N.�-6��4��) ���m w�>^�Ƹ�l���v���U�߽6��B��[���o�vx+=n�Mņ-I����!4y��]*w��%��ߴ��t�Q"�O0��]�Ơ�k>1\Ws�n��Ԍ�f@J��s�9�~f�'��O�10�N��tV��<<�f��T1�A6� ���ߦz�)�ͷu���+Q*r";�R�{����� q��:DR���:�^�B#J��T�&4�7΂h�JqEyL����z�?xDK�D�O�ϙ��`�..�ƷV�7�c�	3Ĭ�0��
|��\k3`�����\^^~�"��Š�?��@��h�M�����7F�aM%�������9ħՋ97��7��pg�f.",����,��2��IhI�	�4��/��qq�x
�D(I՟�J��6?����+l@���NcS1��(ѯ� m#��y��	�mjd�W�o@h�Ĩ!�����Y��A��;��O�8V�A��kL�7�\a�lH-��%E�*|���������NG�w���,�ô.�mv��k'������>�G�r�J�Qۏ�x�)D�q��P�?z�2r��;(}-o��f�PqM՞cy�f���t�����Io�@|�*�uN^؂f��G�����]6>W7qs���>�6Dhxq]��I}��5���t�Ξ����07�q\���X~���HZ�t��(�K��Z���`��l�KAP�5T��+�s���T�:�xbzvV��e�J\:2����%��9����l2����m�ޢ������˕�$�3���@n�D�^e�������6�=q(P��3!����*@�f�ō�j ڃ?����6@k������|[HeM'�����	�sE<����67L�c��W�W>%|��ao�5���	�W۞y
��0�zy}�����dS.ȓ�����{oۆ�O���9����sj�Jx�qI�v�x� J������58�-��<�2#o��qG)��f>˄���Co�y�����Ԏ8�D$A�$�p}��c�Ld^�����Q�d�zl{�KS׻��B�x9.P���CK�O�p��e=�
hii��1`��C��k��|?���[ڕ�rd����I���z���ǽ�����b^
p{m����X�秘&Em��n�h�g�
�5կ������`�_I�vֈ���~l�[A𿭴���?t��lM�S���V���lP��|�7�ˤ�O���w��f��]<N�8Vs ���c���K�&J��<cR�oE�6,ۨjh�1��z���h���s%�gT_�7\c�{\}F�A�r�G�¢Ʃ��3`�7Q�j)K���-ŉ2C�_�ņ��!����:T�L���p���M�ZO[���K���uc���q�%o��m��&%G6�O�}tۈ�ݏ]�f M��I��]�Ҟެ|e]j&�@�T�Bk`%�:�ߏ����ڱL��ek���M%M�?����9�?�ք�)`K�{=B󲚷��`gVUo����7��v�RXu���u�
>���?a��#"#3��\����<y�
��&����'_���/�ݫ�N0K�r��ERl�����ny���r%=4:Ph�wx>�@��a0h��?N�[.��6��x�-�Ƅ~'�j����x��+ڕ�4���="�"���GK@�{�LY��S,C��3�[Y�~iF��˃���1�4��9�'�)��u��v�S��@��6��Z���6�c2+K�v�ve�x��?��א$���	қţ��V�G�.�p��Si1oGP�շp�*{>���
���3�zM:���o�����={Ҁ�c����[��!�~o��2)p�s��NM��w��R(
e���X�V�&{����Ǯ�Cb����8m�x�ń��ȓ'��ƻGo�����R��0��ߏ����+��&��4��M�K��H��j-ɓ�Q��Cm*���s��-)
R'�b@b��48�F�����T�_��`�},nE���9�Ǆt7Z����`,� I%���ؐ{�NT-��$4�ߜb���f3�4�VQ�8^u�I顚;�kh*�����_�u�����0��m<�eػ�wP~sFW�<�A���F������@�A����3.��?�����~�R";#Ư_�%���ҏ�TL[]���I �?po?��1�P��7}m6jO��4��
���y�*�?rH����<�~ZEh�%�E=甒#��o�7�����Z�~pǻ��R,ft��7�'-߾q���~����l>�VGs��vD������� ��H��H�E����.�/�)+ɡ0@G�������wv'Af��g�?N)v6L䦭�E��Pl;�W��ˎ���ҵ�md$V������љ�̮�vwI��T�?2{�T���T�bnm'��-!�:��o�:�^#�?'���嗥i��M��.3�Ʒcy۷}�`T]D����i��+���IN�$Y*��Ń/ U�h�*��LG��fႮ�1��ؒdU���A&�-�Z3'�*r)Lc�Z�	�=EW��ĩ�+�ȷo}��F�,U�ykN*���ޕ��n�?Z9N?�N䣜)���=Q���B�	+b�Q���_/k�c��*C!��E`<
B1��T�	Obd^�נ�[�p�,lgHk����"b�mٸJq�{A���qt�_��q1w�n�p��)^�M�z�)�7��^k��δ�W T���z�LK���}��#^'(%�?E��9duއ+HJ�F=@���ꊓ5DJ
���h����)�z�$y|�*�e�X�#Dp�۸^�+A�\)-�����'H=\"]�]ț\�.����1!���[(ھ�ի�A��˾F��Q�P|G�(�N|�B�U��/�f	Y鉾�v�'�i1��'�wi�>BuM5ԜD�.�󬂂�s��<�1X�-���(?�cm*j1�~�T��4�����9U�E�ͱ47���7z��X�GD�<X냣K�[ɨ�'���20�[�0�p"�T#�9$p�P���W�BI/j^ɿ�� x)B�>Vd���d=�g�5�W��z�9���M�[I�J�y�\�"�.)D��]�J_R&�1\+ �/Ja׾s$�<�7����3zJ1����?�+!�
��2����{'�:VtmmǨ�yǑ�,��,�f�_�W*��p�Q�F��.���`�bi�#�==��+��ٷ���!��������.�,'�X---��V�3���Y�t�J��� �42�ɑ�d�RiY3�*��v��ߺe���_�����E/s������c�i�*��_F~�2F�'�F�/���tT���(�U��-C��jD� zJ� <�g:�'�j1 w��

�3��ZL��.�ߊM�ޒf��򼛑�읝�����y8�pcy���`�j[�|�⊆�L�\�$�e�XA��iP&��7I������cp��j���9	��` z�RG#ҹ٠Lq7~�j3,�U<z�
i��׼����6����3RrT�N+�?��PYD��%���2�<�JD�娻$���u���k�i��U���X��E������Z"�ѳH��~߷Jn���}�7�K��Ɩt��W'Ԁz�XY�/�|������"�v���t6ʛx);`O��7�<�M��70)�<�Ǳ��i���)��U������" ��oآ+�'��e1���x�eNs�JѲ@�ȅ��b�-���OĘN��I�;_��a�V*3  � 8�w���`�3J)�VPP%�ӈ->h8v�J�^ �����v�M��������N����UC�[����bY�>(���/�39a(���'���m�8�[�+�_3#,Z�L�2D2|��-� �G�'C�q���Ϛ�:�*s��f�P�РW�`��}
�a�0��hs7�6H}(]��s��\�T$:���h��~�	�������2�ZTm&����o�à�	 �>�T�s�."�f�BȐG����G��/*�\¦�wCJ����Lu)c�c�Z����o��f��	&F �o;�-�����+d�}zl/+�b��:����@�2b��\�C�����
뒵���: ��!GC�\)�S�,�i����yҼ/��wL�U��P�Kd�2`l����rc͘	���~5 �P��`\�_fжau��Ј��d��ܰ)L��5��R�a�5���Zȗ�3��uN���6*����=+W�]e����N�յ�t�W}�!��v��`�)�Ţ�ɮP�h1�[hک��į=&��Ζ��F!H���L�ߝ��� )OݗT�1�JR��nJv����r�WFi�\ju
�@�Qq��.�[�N�%r�:��;�>ˀ[�~{Z�Iw(.�C�^���5:�� ak%3�r(��"I���/���dX���î�x��i�>�+��	�[�S�a�&GV�p �ub�.���a	R/-��!�)���#��()����ً��>��s*��ȏ��A����(�ם�2r�V*ի�xݾA��+��A����պ;�^1�Uב��Q�Hsſ�k꤉������e�o�����rw�[N�>�ƪ�*+C�5bw?���j;{P4���א�[V8�^(f˒"K'ǐ������׹&Sxca�T\<f�v�jMSqXc�6-K�@�Sֲ!�2��;����ʚ�������Emcs8�M.�p�6��e��$ ���5���}���4�������ƥ��{~��}/gF���+��Y]�Qƾ,č��z�t�`�o�nL�']�g�S���}(�d�Q�ӆ�JXhu�����y+�[ҦL z�w�m?��Ʀ&¥/G��:�2��5�>��� ��5Ե�8�w�.Ѯ+3����h�P���6���x(�:�򍫋=ɗ�������xl���w��,r&�3Z�ʋZ��oV�>P�v�`�Ɋ� ���[HXh	�Z��ղ�<���UW��yMW@��ƣ��{tt������G�����?�B�B��R=F�vwVfw����KU�ʖ𬄵�v,�<�S���'�����U�@�&\U��Q�c�#�쩉E���F�nK�=��e��h����DP�J�۔�L��<[����8�_��2�����&�^w�2v��Ql�WK'X�(,kz2��c�����;��yi2�O���S5�%@�Hխt����1����LSMz��V�x�HZY��%38���C
�{H�'M��@�Ȉ��aӁ>�_n�J6Uq#TmP)�,�oʍrW�G ��k�	�_����n����`�[]�B_�R(KKo޾� ����U�	n��{E����5�_|{�1ѵc���θ�kr�)����wWԜܛ�j������X�%�nK�n�;�
���1C]�FIǀ������u`���uTl/��+��KU*Y��d�����a������ttz�� �M�� ��õ
r��k	(���7^�������A�@�x()���ڼ,���ЬJ�?Tj�d|*����~�L�lmD�$���Z`�Y�ĭ��	9nU�Lc��:g���$Պ�"u�ǖY$�b�20��+��su8�9�ZwU�ɤ���hE~$�į��-�uoce~9�.i�!�������P&~�"��p��g�%<��t��Pc��9v�\��HG��W�r7m-�Z���D�T��ۚ����D��^��M[��f��G������/l�WgUصmBB�;���P�A��k�.���n�ZAbhf�o�����q�?��!�����:��^[�7��	��J(q��䊢�4�cW�$՝\\`�/&6�&Qh�%%'+�tttX��*�<���2i��^l�\���*�m2g�M��Ȩ'���Yޖ�%���t�ѷPuIe�XՉl�oV�zu�R�0r����XR���ňp|,5��.؏o����6NM��U��D�o~���h��0=#�*�PV_yL����e��o���^�q�/^`q����>�˞�
VPɦ�����YU[��Ҷ�9�_��=����o�)�F��ce�G�-՟�����n��羝*F���\B�e-��5� ^��M.�[��|��b�oK�!S�J�h������� Q����߳"���)z�ͪ��q�������wҰ���~�%�x2���߇h�v���c�-CS�����F^D�F�������ۆ�0�`��	ϭ)$[���P��r$��.����I�-i4�k���d���i2��$�p�XJ���i���^���]U���M_pu��vN�'�9��M�O��8��c��(Q|�(''fD�'�l;1�u�ip�eCO9�g~��qSz�||#�8�D<�[ڪW^A���w>��C��Ӻ�HB���|jA��k�Ӧ��>�0P�a��Os����\LJ�y�����?�Ü�sR��^���H��!��U2��׍e�F�?�Jy�������n04�I����L����c�`g³�MW�_�z���6����r!_��][j���B�\~a�B<Y�L>�N�&Nda&v�^��G���xO���	��2���d~�>qV���8d�ָ����d����R;U�s���6�j8��L�՗�1(
hT��
���Q�&��EQؗ�O�Ơ���	���"^R����>�׷���/�Y�ͷ]����P�����N�i롞��&\/#ͤmoZ\�JZ�%��b��+���	�@�+��4-l|��ӓ�)�����Ԅݷ��s���aEߝv/_��oL����]_��C���(2e�.��8E�+xw~>�x���KDE�p�����i~�Ȱ����al�!'��E�a��wwJ�Ȋ���Q��W�B2�M�MǤN^F����܋��t���#4QY1��
����YDu9�Q���1J#�H��J��i����g�3�B�[W�����3H����RԼ����Pb�9���s�'`�c|�F�\�;����\/�<Ge���j���uW�Sĵ��L"���;=�rE�g� 
q.7F�����d�������������˷������Հ�:��Ʈ��j��y�c���$��`��0?�G�h�v�֞�"���.�O��q��;Y(��L�05�@.�~'�JHJ�Z�ߧ&>&�_+IvlqČ���������9������'�5L�e��ni.~�n9����f6J�,ٽP�f.���;N �B-`A�voX(�����сXIC-�U+tˬ'3*�fi���<!"�S,�u����NɬRA�3i0���]���>T��m��ā\K����F�}6{):��,uLuͤ�?M��,�z���z�j�4cS|�Sgթ1�Z����6���ί/F�s�%��|@9����W<�7����ˢ���m�-�[��S���,w�=��<�����k	!�bϮ��|�7�Q�� "��a��]��lB�W�����2ߖ�{�+��b N�uǲ��Wahh6�я��j��=����WE�OkTB�L?4Ӌ��y&��lt���>��ل线�J�AS?��<r	=VT��+io(� "^�|�,�E�
��@ӲPb�9���`z*z&����?��6��5�y��/l����w��	kW��W��+��Xw΃�v[��C��T�2ﱈ=#��M�������m#��ʯ���e6�9������ ��;�d�2���M�B�i��ү���P��-;�F"C
��ƛ4ލb^m5�&���u203���#f�ف���lA�Q9&}L�>��CYg��X�̿�D�M���C�L��������Fç�L�����,�������^�e���m|��Q����ǥ��X�Q�lZ�PQ����ݞO��-ߥE�A�?�Xˀ�� �y�ݥ#��b����RZzO1�(���2jǈ�w�r�_5!3a����B҇��^"]@��K�u����&�"���'�.��=b��y9*]��*1鸫��6U�hS<�{��|�yʖ]^Y�U���)1�n�O�S(�W�I ���ya��E�0����Lb1�/_jHUԪ�+�	v*� S���2K�S��D�/�s
)l�A�rL4�3�ğ�K8췘WnVB��<����1T��sl��%5`f���W\�K>g����v����?7����>�n��7��@b��(m\�\��OO�;T��
�g.�'��2����Z3A��	91��i��${̪�� �������
�����:�qu;+�CK9j�a#����=�ڟ^v��^�ٲ�?����l�Ƿ����
�Eg�=ߏ�k�J�����>.�u�����O2Ś�K��~�#N�O�K�"��+�?� �W߿I��:�5bM���1G���C�n�%��o�1*��\_�I (]�ӊ_��%������X�f}/��ǖ�ءq�ψIH�ShK�z\D�GO�ֻ5���m
���7���V��	������C-ӓ���E��y�[K������5~Q}�2�pf&�u�f֖�TP{?=%䊣:!U�i2ட�X�_�!j-W�h���_-`4�Eh�[�YX�	)��+bb�'���Մ����5�߸X��B��g���/�ɔ�9ǯ:��9�(W���䷋/�Ԑ0��e��f-�r/�ͬ���K)&W�/�ǄU�L����]�g��j�ԏ�~ CU���|RZ�h3}$Bg�/f�tE��Jp��|�/t9��ψ#�vŨ���y�ǈ���E�:)��/F]S�@����J�&�m��n��x�_L�l��E��4��.��[ ���I�:���������So���n�F���r�M��ڪ����<}r����d\/$�E��Qթ�����q\������P�q���>�2��p�ö��ԘOU�Z3f.�gM��ȷ��e{M4�;i%�@�����9�n�Rw��Z���v���k��!�]�y�v_@�J��]]N)o����+�zm�������'��������{�M�Rn��Gb�����w���['���B
�a����2B���lc���:����5Hjk���Dj���K���,�
�g��D˱�M��?,���b` �o�_����>���^E�LÍ�����u�[�k�@�&��۶����+�{,�'�0��#+����5)��o�EZ||"~D�_����p�^��RN�&x6�V��j� )���/b�D�c��
����?��+;'��� �쌂�d=��%������,��G
"��톱3#���CV�hHE��Ix|: �$(U7j��,��ኀ�����$"}�}9��M6L���ӯ�2��ΏHd�,�x:���=s�#��>���5�M��Ɨc��i��Z�?G��f���W�d3��h1}(Y�E-_� MQu��t'�Ʌ�1#�(���V����v ����58O�O�&�b���[� @��ت;�E�;�ȟ��֌�$��a$�*-�Zƌd�8��V���8]�������4�ƣ�1x;t��$G�KG�)�
� �A*��΁����3H9�������ɝ=�����q���r����0���5lܛ�|Ȉ���=^��x��J�	�l��]J��P��hE�L�d4mR��z<���S��76��f~�)�mw�l��t8OZnv�9�;�o#VB�P����mt=�B3{7�@�����5�C�@�/c?2GF�wp�R�4J��{ʀ�j�NU�6�C��PNֿ�_h"��xK��ϣj�Jh+*�˲�ĺx��@�ڊ~8s����Z�q�*<�k	m�T��蕑��|c+�(j�2s�7��kW�.FL��PaYuQqӇ�e;�C V�MIt"���n����P���P�1 Q�f����0}�����G��"�̲��2wq�C?~��:��q��V��9ʢ!N�P�O�*}H8��c��l�J��M����v�� z�g�ԉ�:\ǃ�N��sr�M[��xkn� ��ڶ�C�u�e�lA#��ʵ"�Ը�uS$����g�%�9�ow�q⻝9Y���}VU�z��q�H�i����
�b�
1$c�K�AΆ������9����սj�7�,\���]-�'K7.-F��#�T�|C� /0��EzD�T3;�y�}��;U�����8 I��-?�jh���%(�^��01��I��F~Q�(�C��!��m}�d������D��Ů|i^�)F�C� �����
\��L�Q����0;����đ�|9H�=��\,�yo5�5����F{��dTҶW�����P�Ծ�(�Y���;Zc.zB?照���
|\v�qH�W՗�1����y��t��W�������C�Ω���A&�G�`I������_��F\;��j�G�[�x	���	K����r�ZT^N�l�Iw}������^~cÚ�u��cvܓ��=��R�'��TJ��\�S<���&���<�gm�!��f�$E:���b�ٳ��٨PǬ�όe쾫Xv)����*ѵ��w1���E&}�������G���w�{�7&�Z�g;�FK��t���J��{����_�8�,�+�����(5#.is�6����ҋ>8� �i�V�G�z��.�N�#]�G��x�^-����y�X���ص?����%�&b�65�l���I��8n@I+$%%�DL����p��erG����|ZàG�]��[��!4���T=�377O�������`��+�~K �O�D�HIJX;�b�,K��MN�Wn���	�P����#�ߧ�Y^��p����{<	`)��hg����Mx&4�����u�Mb�M�DW<�����Q��>B~UĘT<�)�l�&���e���^�RBN\K�>F~kD�K��WG���ɾh���k ƣE\>+a��	b����y�x��in5ޠ�=+�Ht�v~.��;���D骽*��W�����m�}��u�K{�Ɏډ��kû��8��l��ޯ�s;;��Il'y��<�Ċ?�4hQch�9�uA=_�j�}ˢ<�$#J��I�E�k�S�&0b7����29n�p�G��O��Xuo��X�'Z!�!槣X�aej
qIK|�a(=�~�M&�	�r�8��Y%O��ڢ��7��]>�*㕂���~��bh�==4���#3�~�;������_7���g��.Ae���#)9�$W-���7�P�>����Kq'b��P{��^΢E��؎� �V��s<���i"�W)�ɲ���$k��O���!� �j��^-��HȎڣ���ȶ7�RH����5�%�(N$�m�I���ӛ��U�����hA	�G��V���, ���Kt�����p��wq@�yD�#�9����N���VA�ۮ�^6�dh0?�l����vxXeS���Jǣr�l{_x�����:���_�3�9<�+O������r#/t�\�.��6m�B�2�Zq��~��L������q�����W�Fu�[�E:����v��y2^�\���k� ����hw#q��`�^�)��e��9�ˑ�
6E�'�mOx�]����%�V]o�����b�id��0||�z�cy ���^|{:\�h'�m�R�M�c\�?d'jF�od�ą�gA���ܲ��{\���e� ~N�j�B�}��Q�����!�ݿ����,l��{&�Σwʭ]ߪ�"aYy�Z���ҏ��W�}�i3�]2grEhe+0Ǵ����	�����;�9���x�_����T�I�7ƞԠ�}9!��ɬ|}1��&4ދ�~B��f*K��r�A��������Q毳~Ǽ���`ܩʢ7��¹�)�_�Z�d��L�~�9�)^S���K0�><���� Cl%-�I����3��|TT��~�p��q�1�sЦ����J�݇�gV��L�pSj�/�$�d�tcky��I��2#��&��0/�LV��$'_�/c��to��K/������s��£����.�T��=��:�;V\���.�E��"��a5��l��G���>�
<�94��gZ/� �%�RZQTR���_��뒯ҵ��Z��S���8�/a��<w����ci� ?s��X�3�`Ŗ.\N��08{�?7��OV��d�k�&)R�y*^��_�딵�)�7(��!b<��ZkRF�^�H��,J�M]���&�"��lxʏo������N�X�t���C��&����:�Ϳ!�x*a�8�f���b��A��LבP�"�J ����Π�z&%9ެa������8��HS�TtSRY��$~˰@�q���Z��KK���IВ!��;��M�g+�NH��609.J8�q�r<����ỽ���3?�i�mrA�9_��rŸ6�6b9�W�g@�$
;�-n)&�n��ٳ?RJ� $�gt��aU�T�k̄��|L�UQ��-����"U�v�v��:���Sd�zfb�
t��:���h��$��u*��O�+�\I�B�����������5~v�!dP<�I�7}�͆hD����$��f�n���w 	0���b3�n�ޱ�__""�b�⡦F�a��ؘu]O���1�G�v���_�9��i�b�����`yj��86B2�+!���wM����,L�7��;��o՘M������1���^�2>f�ѯ��>]���+�^7?'�lg��/�5��C�z(3�l���0T
�2�
���/���;\�9�&}�g��p��&�$ZM�6Y�B��
��73��!��ĝu�o��F��
����Bkɷ�?�v_e������|%j���� �\'���tMR�+[?����� �k	y�ʩ�V��MW��ƭ�BBT�e~?!��r�e;�@0p*د,:Iky1���v�XJTN��Kb�O ��;K�`�2�L4@j�d��]W���ְ��"��}��ރFlb�?:��yx�{.�Ø#n��ˮ��Q���b����>r+���}艌��sRw�0�F���a���>�����τ�Xk��yV+nV3U�KdG�3	����0ΟnW4tX�1;�M��B�����Q���O�Q��0 U�������02�/�l�?(r5�pwj6�cμq��� (�;�s�%�ς��P����� ���[��v������7����%o�ɹ���jH�1:&����B�˵�ը��4p���v �D��n�]�o�H�$�����[��f,2DnFN��mBn�,���r�ÛP��p#}l���O�@�!K7��撯�#�ڲ(�x�-���=��ac�w����e���������� (&Q�����:x��������Ä��W�q���j�3��u^&pɫ�F�Wbs8D+]c��|[�����{j�h>�6� τPpڌ���_ݤ��5�%oC����S�	�Y�M�3�D[��np���x���iU�)���XH�콶�����;E�au:�t����G�Z������4.s�?(��9<��_�%s������~��j-�v�hj0��w�>�5`�[�"B�Tc��'��_� K:������?���քi�{|���2P���p��s��Q�7�6��?c�S�V� ��S��i.�5�[���SJ�HHC?��@�1<`�K��bU��D���ט6&߱�;j��"���|�w�v�~��� ���Z���z�㉙4�n��W��j�n��<O��l;��$:��*ĭa�lsu���Ͼ��F��ֺ����v������.�bhR�� [�M*vOr���+l�K���Ӵ>-��?;�<ಂ:.'��W��▻4<G�h�e��Vb~���k����Y�}8��/�O��[߾<mF |����I&њ�h0ӄJ�� �����_�q�+�2?Fn�P���/�=��j� ϗ3563�<�\ILpj=ѫzD/�����^{'>u�#�j�aȏN0�l"����@)����}p��������h7J����v�'#��C��:��|_i㣈�btK��=8�2�d���t�'̔r'�L�1ft�����(��DRm�i����ur�W�'��b�X���[���������.���j�Z��`I���o�iU�K����%"_�ϔt��3p�R�e�v�r¼�]�kT!>����`�N�{�<8 %, D�a�2aI�X�BI�D���U�-â�_��w��%>`��Ä�U�kk5p��Ov;�!#�>c���X��PͲǃc.h����s�
�=�6�	M������
��*��4)�cVR�3D)p��UF�'Mo�Js貧!���"��浒"4A�G(��mIaF�2�q3x)n�z���巛���� ���{�E�LFJ=�HMWD�P�� �)M������X��2'��*�~ђ��E]�_�\��8_I'{�]�{�:%��>�mC"�s[�uog��R�,h�Y��������'���H�~U��S!T�xĘ�w��n8.ܨ�9�z��h!�l_�Z�e�`7m,9y���]�y a
p	��NAR�E��e{~y�DM<�#$WS.K��nY#s������Iw�!��/���j5Y�5��p{\���p�Sͽ��:B ,WWhx�H��Y�QG�������5������]Rq�).Gm����z��=�ԟ���w!���t���~�+�[��w�sd������|����W�?�����W���xqF̈́�����zC��
`�]�+P��[)��o^F��?`��DZH����a�.��#��YLcV��T�.&��~��#P�'s����AX*RG����zZ|Fs�aD�k&Ew��stQWO"�_��y�0W�\�4��,��������$�b�m~���M��T��r���X�Zl)��7����

"6J{{�鴐���5��w�����[,׍��G���n���|H���[��>��ի�&\)0�s�ȵ^-��$��qG�R�=�|��)&G�J�"��ђO��Kӌ��vy`�7�kΓ�Ԭ+��ʻ1�]r��k������1�r��`�&��m.��wc37���.&~��2�Kv�-e��K6�٥@o?���*�駔�W���;}}E�G_����c�첯H|��2~�ڃQ��eV�M9�j�Q���v��ǥF��O�H�=��^T����@�pu�pr���|���0\rİ��
z�UZK���3��~��խ;J��1��	J��0����n��t�.�`�����5��� EęfV��4oꦎM����?<u<���P����'6������ÿ��Y�ʕ��^�>t��D	�1�Ѱ��g���;�{�m�k��i��#w��W�d(�$g�J@1��
����]�ծ?@%4��,����V��������)ߺ�bܰp�R6��'�+���t~06�A����/�����B�B)�P�5�k�JZ�Ӣ�F��"� ?��#�N�O&��lyU��P�^!j"ڧfSV��SS��(6����~}���F�u����&R��}��[�{�^��x�<䖂M�+ |v��z�x�̯�31�V�vA�\&�vR�������^فbm||x��rg�Q8�����{�Ӧp8�yۊ�b,��I(�$ML���'���)��T�<��66�گfqz�zX>����0N�����L�y�z�|ۗ/{��߱�������~͵<w�G���[vF��d���?�N|��}C������ 7R~u8�1�z�<�R���U��`V>_�#��,$�j�%\�i�?4���@*�kR�ű>A �D�r0��{�x�e)����շ�*�V)'�3���ר�MQKTS����^�L�X�>y�!s�p+�&c�B���36�0��x`hO��6ﯗ�(��q$y:�[�{�z�@(S�K�.���j����[��.K�'�ZZ����<ңnÙﰠ.�ǤU�AI_t�v���Z��T�6t�֎�σT�)�y�6�P��Q;�U��M�
����&�B�YG�A�{�����Ej{����A����Ƹ��A��c	����օ�~ �.2���$�1i�v����2I�H�,�ʙ��@m"[��,Y��ul��^U����;��tL�,U�d��	���)���x-�
��.fm&������o�M$�d(Ω��m�c�^R��2l����o}Tj������UT�#�Z_vfO-z����q�c�.��Kws1:����G�l!x�{��=E��L	�!���0�p�$ X}��S��_��S���v��1k��Ӯ����ۑ%&�X�e�{? ��Z��:X����|�g�D��E�g��$��a���^)ke�f�Nֱ��db���O�� F������E�2J��w��|a�b�]�B�{�36�Y���C�sJU3�p4�	������T4K�&�Q:%�e-z����u��W)�	E��|]Ƚ��Ձ���r�sXG\��}괏:�����^ˑ|�LH��Q��kJN���ϯ�p����J�� #n2:ح�qc�����DV�G[�]/�oP�Jtm�����^���`���G�<��sge���o����*���I,y0�B�6�pK��.����>����~�����7o�"�6|�n�?�0I3r_�� W)'�]��-�|ɭ�".���5��J��<�����<�j��L�7������>�o5��5�pӞ)�ӧ�����1}W�j��̞"�,Đ����!r ����#��EU����8���<� �����e�%
̭�h���:T��2�ě>E���Oz]�/�W�j���� �X�ٸ�'���.���g��E���~�H;if��5��.2m��Jv�9�+�%���}�IkG���o��[��� O�f�׽�Zu���f�$,�?WZ���*0Q��+����g@$����mɃ-{�x2�#?��~a�����g�J"fe�d������t�U)UY8c��Y�����K�TB1�����bD���U���v���.�|񁑥�!��@��Zz�,�����S���|Mc�����S�@3h��
�j0λ�R�#�#7���2K{\�\Ӷٛ�S.:̧O�!�G�4��[�
�)� PL���!9w�(ʂ�A�.���b4�y�	1�qyq)=�Y��s�n��J)i�
Ƶ�ٙ�8�,΢`Z���G���s�p$t~.R��]��l�67����XV�^�|<�J3���c��ȱk�q�� ���_<�N���ݕ�h�����|�)%* �^\�{�m�Ai-oB^Bi�4P@9��v_i'�w�����3ʝ�)L�*��r���?���~��
��n����Q���*A* �Z;iP}�t�&!���1ޅ���U���DThd!��u9L��^�Mx�#4A��0������Ur	8���;)���[hp��[�Z�	���i�"��3_�8��QJFJ��F�����5��{t>RŊ&�k%%�xQ�'_} �I�Uj��U��Չ���z2pe�Zu��ގx��!Yʘ��pEf�,��
"�d�wE;X�ʄ��6�c��ɘ�����l�1�O&�v�dP����l��O����r�ǥS����k,<P�f��g  �"�<O���mN�F`��`��,���A�
C�4�3:��*���pSA�[P;Ƒ�%��Y��_i����穾��Q ��h��<�燵�5p�/����)c�J�7��V̎t���j��r�1&r(e�+����L� ��};���p$�LU���B'�x�Z{u1����M�1'�O���%�u�����34���|T�,s�Ս�������%B�Z��(���h�,yp�<���?���nE���d)}*8U5p�G[�˚/�ۇ���b������B��L��0C5���B(ʺ�+|���H�i�X�6�d�D�9��U���#&u�q��CF�L׼�����F�K/kJ�W��I����N����=n諷�$��)�a?�0�z�/�S�X.J�ѵpz}|�[H�	��X���Ñ����'u�-� �[����T�5���{Bxl�K�2A��~[(R��i�D���b�E�4�����cC�D0~�G�ۜw�/������9b�8�?jS��՝B���ecmR+��L�ɭB����-J~�ϟ�Z��x(�yV����*��s�@s<Yɩr$Ѩu��I�@�اgt�c��aQ����1� ��+�>�wN* ���+�%�Q�D����ҁL����P@IȲ�ʵ{��ٍc���^��>x��J\���m�d���pNM�p��b��nqujꝩ�>��w'Êj���@�1��7�O" ��ʤ!D����)���������-u O{�Nvծy�?Q��P����<����1����v-ܶΗ�9�.�Y�������FO�d�_�U���JZ Tj�yV�@υ6@Bnؘ�v��վ����*���ь~-���*�j�����["�ݥdb��;����N�N�����v��1c�B��Vd�#�ls.��f�H�=����������)3s�� @��6.����T|�K�>���Ю���o�'��a��z�SM��j%�l��%�o�8���%���
���zٱ�r��c~�4$u �U��i�+]�����b��L$���������C W�p[��P����O�p�ؤ4�y��'����$dd��M��v��x���:W��v�����:D�Y��(��P����t��U�����iR�g�»+Qw*��%G�q2�q)!��}�W�.�����7��78�3l�6S�ȅc�L�Gߐ��֍8�^��C�K����w�Y�
�}Z7�F`D��ش�?��a�I8C�G9�g�n��"�6t�ԖRv+U���������%�Va�i��᧯þ��?5Z�u�t`k��Xyyf�t�y��Kpf��Ң�;�>�<����Q�8�{|"p^�����"�yM&v���iz&���3j�7�S��5ISZ��ƒ�N6n�	�t�2�:�Vg�*����V�<LB��roB�d���[/7�gJ;I�&��3鰀�	����-^���4�Hs��*�D����l`Bj��#�O���9�6:x�$Q�2�����Z�ּ+h�!O�~>�+���ͳ���ŝ��!WtI��)!��6�[�,����Bv#ؔι<=F�#"p�NĚ�� �a_�qw�;���=ɪ������2릚�ʲ9��ƋAmG��,��m!j؄���'4�E�8��GAd�:��&C`��߷E	����c��?��nO$�'&7����L��hhi�}�(�΀i�z�O�N���PN�ҤY�I�� �C�d$.B�b�s��9�*ي�<k��}���p�U6��1c��/o�%mT�3��e�!�g�_Ci�˩L��}&���(15�����4W��,$V�������&I�𿠪�3Q:��d�~�Bsk:[�?�f�R�Q�4��=�����ۢA�)at��`\Gye����O!?gȫ�>��_7� �o���ˢ ��|1Dߋ5oB���B5Ip.f�'���Z��i����k�X)����7���̿� fn{n?K��K@f��W[9G�$^�8N���
RhU�2�0-�
j軇q��s�Ny��0�X�y���N��Q�4��H��	�#|�7�)Z	�Ӏ�L�����!�54m�F�j�[!}зi����љ��f����?���?W��s��4�5�#vu?��u��z,N�y6����=V��bB���"Q�瘵|�[O��h���m(��У�9��o�� _*�u��H�k;��vq�y�N�q�֩aL�"��]�Gγ�'��\�5����`?��R]���\N�$�������4��s�6X��.��!ܝpU֗\��$V���o�,5��2v��i�r2<I\�\�e��1��i ��d��O��ɜE�>��||�H��֐�T��#p�_`?�J��5��jt�&����>��o���� ��p�J�W<���}���Xγ�A�N���}�11�в�w1��Y[���D[��I���Ƶ.[�f�������$�s&G:��N���؆��Յy1��b��b䗚��E���m�bzK�r�E܊R��[\/-{��V8�
j�����î15*�Ѫ��L���M�C1_L鰫/das��(@S���p�q&h��-R�wg��.��I>4�x����[�Gzd��N��U�*�%X����B��V�$�.�Dd��r\��GqW!�@xCL��D�5�6#�⡧`6��y�P�?Ɛ+�������d��;��٥�F !�#8�*���g�]Q�F:�J/���N��XIMJ3k�z�A�i�xrYr@�\e�B�7��ߢd�-������z)%�Qg��7	�!p]�	<
Mt�z���En����R3�<�wD���E�����w&O�Fk�Sԙo��<������ͯ� ���f����g0������Q>��PO�dƮ3N��IG>_m8�� ���xC��	�I�~1�UE�,�'��k��V@6;��uz:H��h�(���s�k�XA}Δ�� �}c���[�!̫���?��NNt������� v�:,�jXV��0��A�.T�2��r�7�}bx�����)�.ZJ�@]�D�ޯ]b�ֱ7���⦱�!#���)rz�	���7S�td>���)*��#g�ڐ�6���%��A��#!�����{�G`�锛�f�ǧ6ѷ:P.��;iǫ?'�{M:�����!��:"�ʆ6W�ݤ�#�V\Jѐ��>�8�)�vc뾋���oi}l�</�q+�Դ*��=%!��-��ˠ�K�^���l:qr;��t&F_=�������|�KT쫼�)'�����
�ea�� \����5��O��۲t�F�~���:޺��(��!C��-ˣ-sɱ|�볉�*t�Cta�:&rJ[�%�لUiL����8�L����&�"�ML��V����oP��S�X*�N4��l&7}}�����8ܿ}����nT+urm�@t�2�q��c�S�a�;R� ��<�7�$�cC��Q�(��ǈ(�P�t���n�����R�zy�$����������P�<c�I�&7݀�L�B_�
o�6%rt���'�79�eP��  F�5i��2�r�o���Sl�)%�;��K�.=�Zk�4�PGavdHy&��$z�����Q(f�n+�,�_!J���*Y�.������Nٖ���R�|�i���/��>�)����^`����ѵ�j~	��v��iI�m*�F�~��NA����8rD�Y��/C�;�$���H�a(�8��2��k4�@��<�����61����� 8�u
�)[�/؄�A���]�T&��o^��,4�*� �"���z��i��>;�<I�lj"m! A7 �zm#��Y$����`B���ATu4,��|}��'������+���Ė��Ӵ�]��|<a��fC��g���'��K���1<�$=9�.օƚ�k&N�V�w��A�ٰEg�u�L���������Q��S�-*ܚ������x�4��<e��iÃ�ҲJ"7��k�w�]��˽�Z�n�΄��WX���b�J)T��x���9B��2�� �ٱ��P}��9b�x��,�V�x�*���z*������j��6������d@y$צkF�(׆v��4{.��ތ׻(�� ���&��b �����.o�/� 7f�0q���m,G�|�l�Y�u�D��	C��������?gz� #����AF^�>.;R��V6/�✉��r��D�/_�)�	�^T;���,��t�.)���@���ѾFԦq��yu��TS���ݞ��ȟi�%�������5�Gc�y���z���bU�J囌���d3�D�Q'"�II�h�W����r���&�֏0A�"\�t=��\ �����b?&�'��X��}SH����)$�1����_4̹x����z��L�׺�����$�#�E�ݷ��1���j�}P�O��
��3
ܩ_���[�S>61��r�c���s��m((�l˗�V��>Fl/����M��?�Sydp������1ڊͷ�#v�@��$��&��џ�<ja�����4�����=������4��s3~�r��->Tq4�vauvD�&i�����.��i���c����YK�Ѐ����Bg
�6��t�Qwk�Ŗ���zHs��N���R�����j��o3���l���o�Sm��)@�|��?���a���&D���溤��r}&���Ӻ�Ҷ�3�(o�l�Β��+{|mb�AضH��V�C�w�����ƽ��!��|L���h��w�Vs�ly��~���uHV:����ļ�����Ŀ�OVaf[a��R�0�8mz��3�6�bad*��޳�?�<Y�}r���G�*S�܃�?��t��!��@>;E7��`;�/e)�@2��ׁ'ɷ��qf ����zX1+(��$��dF���?���Mz�j@���15�٨��\b��,l_I�Q&;��%g�L��d0^�{��O<�*����z��&���V���
R($7X�>��ʓ�V�ќ��� ���d)��.^F�8��/�V���Yge��{J:��Ci@:��F@�[��������N�������|�y�Y����������{��#V����04n������hUU�g�k(t�{1���ܴ����R��������Mn�b���,�����g����:\���(��`����R��?h{�H	���q��ȁC����|gF�鲗�B(@�A��/�����/��c�l:tl�r�j�&�x;0 y,q�Q��z�64/;�P�Z�T�J���?���q-����:2�r��X޾�0ܟ��`�]4�O4�F­�Q�l���L��.P9?�C����o�X���a�ט?�m�o����.R;D=�~�M�@]�h���K�����YW��l����ʝ��"ZO�4Y��� ��e��P�J� q�ן♹`Z��l��ՓO0���fݰ��?�����ֻ�<u�H�P��O'�viM��C@�M>fq=�,�b�tƛ�!j�-#T|�m�� ĜA��6��12�`_���˽�����d�%&���ޫcN�ZMG�y����s�`�����I{��>>.j �t���n@~�����
�����@j�lC��G+.��s)�N�&�a����i�s��X��e�_�ȧ�5���VI;�W/$��ɭДWniAV���d�B[?R!��!���70$|����u�06����-E��`D�u�֨��G���Y>.<\�98�l����mk�t��9�Oߤ*�#K
�ɏ���Rp������m��gR���[��̽��j0������X�|GqZ9��똳�:V�g6WӜG��O�c�]�Ted��<ԟ��p��-^w3���m#.�(��6�]/Yiԛ�&��v�n�Js����npl�q��#^b�0�Yɵ��s�_�ٯ��b���r�ΪZG�v�B�i�̝�.� �)iո��h�h��Lq�c� �ց��J�}32'��W]ES�G�����ԭC�P$�uF�����b��)73�%�����ަ���[�{̬���t�����sj��P,�O�c�[���TUqn��S�f�
/DG��,)Ut�fӝX��=c�Z�{��?'��"�P���=ϗF��U�,�w�'R�S���<r�M�v:b�K��[�z���)tXK�s�ᑇt��'�� ����l�M}��s��!ӯsl�E�	�� ��q5�����1Ti�|��?�-eC�˙��z��n�U#���J�j�7b�\R�����n�B��E�����:�&�qMM�7��+ǟ�h[~����l�|���ŭ��?_i�D�~5���N���:�滕����m`��uƈ����|
����Jͧ�(�ףOs_�,�o��Ln6H�۪F%��D+}�Db�Y)Z!_��++��~C�!>���zO�r�[��k��&����3ܹ��8�q�ד>m�P"K^�+��\g���.��H�kw����m]]c1
?zu��E�/1�q�;���n4�C�lM>�Y��hoY��9R���-��ZU�ۅm
�\�I:%�=�}��a��U��`�^�ޮ!�5���B�֝����G��1ű�3Ѝ��,�>H��c	W�=-#B)�Zv�V�j��w/@�;�Jr
�O#'��-��>���
�*��:�J�Z{��N㫬�ۡ�(�x�m-C�^
j#kz��^?[PO@�pG\U.�^)1^x׋�Ef�\�i|	�����qad�	q+{q�]וrh��׎?�n_�&����Y�g�_��eh�C����|LW��ٷĘ,p��FW^2O��j��^���3T��^�Ѽ,�6A��$Om(h�1�]���~|�X!wG�kt�K�%�/7���~�ڄ�v;1�Y�IFI�f��vG���gBG��7O|�ƙ�%���.�N�Mݜ��ȅ����ѡ0���E��9���Q,�c�pk�pB�+]�p�f˷�1)����aa-̞��m���N��j�zQ?�����U�ʄ$�=v1���aP���>i���~��2]����!Fݘ�ҵ�
,����[�����.`���g�c�y�]'nC���%/�s��ď��t��'¶/��K�����a�N����t����2Hx��d���VX�`�o�qA���NU�oCBH����e�����������;-o�\��
��|4��ek����Rbl2z��7�e�l���Rmv������n�6ٷL,��?yq��ի&��q�d��S��}�hS������w��M�`�M5)���u����rU���}w��AT�x�%B�}e[��Q�J�M�o�� "��3�m��=���[�d�0���sf͌1��E����I#�� �c�i�/uhI�j��}�ש���_���R�WX(�ٌzw�|��8������<<e���;^�����F흜|=L���f\jet�9�W]��3�=8�Z�����}�������H?�&�Q����d�M#��ݴ45�+hU����ߗ�|w"��t�r~�Я�����*6��q����S�K_�n*��N�]ɤ�ު3a��Z?f�g%�Q%5�^��VD����8C�J�7R����T��F���(�Ԣȃ�iBbx����UB�kcJ}�?T��"= �`[Uu��v8�f[�a[e^8U��z��c�c�b7��1���P�NK>I�4i��V��Mo\��Ȟ�8��+���r�z|!�����E���Qj��o	��aCcc��V�%�[�wJ���yp��|Յρ88T:��]�/%d�+,�%⚍�So�j�?m�+l�����yR�ӂI���F��d���A�H�She�օ^���]d�࿊�s唡��JMF�)�E�*�y��c�VIz�a��[��(>��P����P��O��� �|=<<���rP�F��'m�$�n��Xi��*d�X1xP��wj��|=X���i'V��>|N&3Z��H�����@6��T�jl��[^�q^�$>�"���|х����Uݞ�U�G�h��J�E�ԓ��:�����5�oK�@g���]�**�F�[�-�˷Ho��uՎx�薬zT�fb������hm~���Z&6ij��U׌�1riX�Wԅk�{`�<� �ܥ�3�>����N1��uL�"��j�Ed;y���EZw^'_�E�l�?�����Bgg��B�n�=�c���۞�C��Ɣ7#�m�(%����Ӿ��o����b�sգw��ʒ�p���f5Q�ɻ9pq���]�-����M��|���S@'�|�κ�T��Ȳ�ަ��$��x>*�7��C��b������� i4 $�m�����'#m 4���Oc�y��T�)����i�{J)Ux��2�B�@\jq���/�f��P�� f�
9�V��֖��XGˊ���Qlr�� [�8����o��ɍp�T�����8~�k]?�t$<OR���&���2��*L�1(R����/ѭK~R���iI����I6]�L�Ϗ.@�=x�J߸�k��C��gwf�v�kd�{˵D�y �xG>�0�Ǚ��Q�^?v7�#�b��3�T�4��*j/����ҰPe�[ �n�EO]�RicK~5xAŦ�p�!���e�gt��X����V\�Q}iB�SJ��^���=���'*���[�_�3�+���yn��ތ�������u��5I�<������a�)kTͲ� ^��}�.�h��O=��d�lz����Pe]16���үsC�FY]�r�ܔ�F������4�ٚ�ܱ�m��j�pβK���\|V��:8ek�O�!�`c��&�v��`��rـ[Bd8wA&�����Դ�	�'��]�EO��/�嵫��]��;u��h�<a�Ẑ׫����x��ߧ͹N�`�thT��~76�J���5�}k��z�b�A���������où��e��%)H���hW+m�յ�r�1��~B�ڀŏC髴fg;�8��6�-�֛�(O3�4G���E�d�9�T�ߍU�I;}���0~Y�!	Qw�5��=#��[�^�e��Y�A�t��������#�Ӹۛu�S��v��t���~2�4��3��P������|u�J9G��q��w�E����ؽ1�v�0$2T��\�B.��x���{q�Ҙ��v�����ڝ	p!�g3�k|m�ϗ�('�)3�����\7��;T��i��Gq����O����@E�ko&�Q�n\}�Q�Ap�J	瀼M��Ο���Z�TM�7���,�)�~�_a]��vB1=k=/��^�z�3�T�-`��������������Ț���LW-t��k]%��,�x
D��w��d�8��] �&��
��IpӘ�Ta仺煟�Z/2�Jp-����+���r���`_�!�m��%�[�$u�Ĩh�BO�����\bo�P#�E	 ���&o�]�\����%���y0�"�r�ằ�~ΐ�X�|Ni�Z�����in���l8US�-������zn1}k�z��|�],���_)גJ����5��F$�C��Xx^ڠ�����d�����r{;Ǐ��Zs3b�O��Hp�V�<����NNG�*�Pﰰ���^���f�?���o�;@����_x_�|)�p����C�s��4I��<��|:	Aԗv�鴈p(���bD�zZ�M_\V#Y��jo���x'JV���܍��Q��i��Z/J�ᨍ��.��
W=B��r�B�r�K�����	��gw/r����wM��*���V�E�˫����^�vŌO�Ӣ��J>��'fʯHr&=�����((w�z'��۽����8�����������N� ���؝e�͹R��^��[�cK@�r�t-jd*ￂ�"�F��Ӟ�\�:���\���l ��T�_�U7ZkV�e-��a7�Ŵ5�s���P��`��&�2�/%�����7�=��<�!��r}.��f��v*b	V��.J�0�q�~�Wb�@�<�`�tW��"wٸ��.�����b ���v�����s��n����%U����*2>���a{?�Z*ҟ�� �A>�H4hZ��d���Z�1ĭ��o�)���-��Q�_��)����up�E�� 
~�� �`e_��������I#��HQT����� �Gч�8��/>  h&g5�$����])y>|�O5��1��24�[�RGH���ǡ�?��q�G�205�=�C?�m=hb�m	� R�/ a�o��}��4�=��AfJ�{���:H�OW�kz	���g���##��f�BKE?�X��G,�BO�F务�C�n��@�rE�?����}�dXq��IYX��Rd^�SG��
��{���M��R�N��Al���>u��B�q�<�@d�\���Ɨ���g�r�Fpn�Sbi >��Rg������;�zj. �g{�m�J��Ӭ�#z��Bl��f5]�� �p
t�t
�'��V�(�ù}��4�r�Dw�/��˯��=mg
C������� {%��\D��[�K2�㋐_'s�e��s�K��&��?�x��*�L6�����mq鎓��H��,�G����o�8�d|�w����K<�,�fm:=�R�&ޘr��w��ɀp����¡$�޹��w��<�J_s�]��e�Ž=�uT��:�vO�'�ic ��K`d�g��ȿ��r�}���♫eT�����O��Kd�Y�����sk�~��`k�D�f�@��n��&���������`����|e�g�\�%�ˢ���,�Sl4_蜖���r�9�_M5PsŽĉ]�+��9M��23��qQ����r���w�a�B�;�b���� ]1W&�v!��h�LQ�w$n�t����Ӈ2���������D�UN����l�H��u3����?�P.�}��j���QSX
C��Q;��*�}�����ڃz�{I������V7��=t*���H�X*8ɚ�n�D�'� ��a�c��pv�N9�B���+�j������k\c���0�E~�C��OL����.a���N'��ԉ!�d����Q-o���/�ݜ߾zN�˷�;N_I��\]5���MR<�YRA��k䬯��tˍ\x�!=�5/rG ����~{=e����ww�E� ps9�4��\��M�z:���V�~,"#̧��#�F�V��˵ٰ���A��=C�P'�7��[]g�{k�Z�Ҋj��؏�<�^���(��I��/I'\���P�c.J���	��~�X�Fˁ�v{��U:�]�����|�f�6��u����}Q��	`��iWm,�;�F�W޵�����{�q��7�%��6.�_��1s%	���Ү�y��t´�CR���,W��U����=�4��\����C��k4�)� �
1�D\|V�n� w�2\X$���+��Ɨ��fK�����ys�4��m枪Q��>�G��D�����c�JzK�����;���p�QC��
��[��_�iF�dk�'����7Vo�O��n��oVA�W D��h�@R��O�N[��TR���{�a���6N��'�N/�Z?�c:� cdt�����\]t�6��������̯�����Pj�hCM�478"0�(Ӭ�P�6GL�2�f6z"j�J�z/�[�"�@7]�+��!!xa ��-��q=��z���y�|���ʀ����j��1P�|��ɞ/�b3^3�y��%A�p����^�Nk�G������rAwMtJ��P�Z�#�4��{o��m��ݐS��P�Z�X#���ؒ�����*ҏ�vd������6Դ��v~p[B+���zLi�?��K	�9�x�{XoB�釬.�V�m�?A���֪]O��d���v:#�n�$�


���9�}B����'�>�oOo��z��/�,i�_�fD���1\9eĠ����fx�]�}�3�A��,%�°�	+w�?�N<r��h�����$jۃ|~-��zۂ�%�Ʊsi�XC�z7?�����'����՟r��Pd3�^��L+Y1�/�s�bδ<�X�İ�+����z�js�P,e��*�/Q�c��'{"O7��X���W)�K��n`sA���m��	%������T�[A�ˀSZ�m�VX�u�4����X�����(���1�]xe)���Td���泉�f���'\�y���%�_�7f�
3��D��h�k���PОf���3F���/�U��A����9���2�n���c��F��wL|@[��-�����x��R^!��h��x�/^���� .C��A}\s�=�ex~&����̔��M��_�_z�V�{h�F�4��<� �E���9�[�Z��QY�\��%��@��C���<�kJT+�z�;���I��&�K�j<7^0�}���X1|�+�v��D�>sϏ�����<��1vu��kGBQK>�G��JU��0�<
[��`�X[PO{k�˃5~78�+�eY�+�6+�gK��<��|�z�4�ƴQ���#T�#q��L��m�çY��|�{�̿}�Y���G�0��*5WQ<���������Ѝ�����jݢ�"�G!�_Dhř�(�oi����]Nq��j��6�iy�`�V�������	~�/�����_�������0\�4�"�.�-�&�t,N��sK#W�Hx�^66s�/N����`K*�?Q�����z��6w��i��l0��� 2�@f)����1���Г�3�ni
3:,�#]�gB`�O 	� T�~z�~g�7�*Oӣ����6p�ШuC�f ����{����%I#7OjZ>�I
��%��l�6B��j��F���E����y��
�$ckcKj��W� mӹ�/�2?mivNƛ<���L v޲�S�u��"�jr�7&�bS�g�U�0Rw���ђ��y�˷�:7K��*��ؓ�!T'�$��O���G�^�?�7�t]%l�b���:��aDĝ]U-�~��eT�8ǏA�Hἳ�P�����ge�����kƸ��/� L��s�<�}	�i��K�����.u��R����(��@��*
�[�}S�P�X��ea��n˻�� �G���t�z=0禟Z���8&�&�ψ[7�`';�{&XX�9�ּ8��l�� P|�6�%���G�����Z����q�6��3B؉��P�rɅ��f�7�w+$�N��G��"��^��V��)�Lݸ�8��}C!]�P ��ՠ0I��w�rT��K%�#��[X?ԉY�Pa	z��k���N��<m�>�:���˓���m����A�#�.4�8;���X@x����.�]�ޜ��~�I]::&!��X�P����l9c?����;Տ��[�]؈��yeb�$���f��iwf�p*����$׵���E����K�`�é�Rı�q���%;��rԸ�/�ݙ�1�:��0��y��+86�`B7w�W���16f�.o���kw{vxuČn&�m����Qs���0����������}M5�h]��|E����K�1��؏�!�AS+�G:S��9��cG��zI�n|�ni!{���m��_c���L;t���@������>����T)�*�1���L��2��/r�W�f`Q7���Q('Ug�g�i��l���<02�3?�l�+^\}[��^y�#�����R����ߑc�ti��OFU<���#I�=b�[I舲����y)�IW�"�
���� ������?8��^�E�=�U4�����g=�m^��'�Qq���G�'"Iv�6"��kަ�n��%<��U�G��2���Z�N�Dk���Z��֩&�[� IW���b���
�%A�E�����|]���I�����"�����X��s\O�]&$���߬���E�Ta�l�*�I/�2d>.�s���NhwS���)���r	�##�z�Ñ�)`���X�	�_T(�$�g���Y[A@�2\����s��Q_u�/��\/�y�'"v��	�~�o;{��wϸ�5��]�U|MHBԿ��C=��U.\;L����[�J�y#VĽ@�dJ��vk�y�"���U�� �<��A�YHWY-g���L���ij��t��s���>F��&�ҁ�(˧������?|�������Ps����;���ݼ�5f�����m�$
Iu�QցJ/�6]��o���In>�t=J�z�_}t��j��- /Yy��6���v)�Y���x{������)	'��}1 +>��1����(�WU�Y��&�d5E�dҭ������ߍv��yhW�g5��ѯ�������on��0��3uqKߥ}��Puv�y�-����V=z
�7��B���+��j��"M4��<�u7fUY�O����ٍO��$z�= v����}�8*�>�J'$Ff� ��q��w[����%Sۚ>�_9���4��.�O�R┶���𺧷�(�����=Ր��^�ʨd������.���2�5��h�p�]� j�����v<2��J��mb��^É�ä��$/�P�����4�z�K�@����K�_��f���Y��8z�zGY�g��;��s�Ŕɓ�z���j��l8�ݵ��u�FI�E��ZR!k�}��8�[e�5�R���[�����1�f���)�U�����Y��/�c�~P{}��&	$>w�u�q��-�k�����*�4SB��%�XSQS3,11���e�\T#�+�m��(,�Z"ngW�����x���n(ڈ�����+��e]D++.,�0�O�
r���#��1I�cccc��K���� ���|{��osU�v��X߭�c�S_�}���e�u@[�����U3�(=�"ޅ�e��X��Je΄v���J禨�����TN"�n�(0U{C�{��FؿN�
1�� �.�A�X���[^7��G�Ad�iYp�)I��}��h^��v5a�8SgZD����h�i$~Y�o Y��Z�sюb���t�Z������-kV�d'�%0�DìAk�9/f�e�U��fƓ�=&=��-2��ZH�?���)Qʿ?�/��5x� ��AT�Ȋ$�p������	9n�t�.�%oFi�} 1�	L[��[N��׻K��o}�NIţ�B�;�[����گ�-��c�6|�F��K^=�'8N`	�Z5f�qa���F������)���{7��5���&`I�J�V܁��]�ڑ��v�=��@�V��Z�6��y ���������������p[��ꠧ�(��]������I�@�{'靖
���(��"B�[=���"U��{$��$���@JQ:Z�Gѓ�CKMK��L_[:F����{�Ӈle���)��i�Կ�?�]����qѥ�s>lro���!�KY/6ݭ�+�uکڪ�<�L���1Ϲ9�fۺd[�;[�]�Kv�Ԯ�++}��wM���v1w�aƭD13-���X5�_�3�D�{�fh�b�EYF����x�8��s�Js@��f%3���X�=��+]���(�x�&�J�UT
���e8h�v��99I	6��j[_�Y.���5�lↀ�׌S��Ef���o7O7� bN,nU�������]۶����������nY�ڌr}4 ��\��S󱝁xH� 6������<2��H ���������x0�/A�_`���UzRRpz:����S���l�b���RyG���]�Tja�4��u�u��_vd�~�����T����(�r��k��P�;@�7��Q�D �\�pJXF0���5v���-���1x�f�~b�|�S
Ձ���=����3X�_�V��;���D�Ypɪ�(�	H�Ď��/p� Ң�=�̰�bZ㋯*�"Ű��g�,�����|ݮOxY�1���6�3��D�F#�xSi��ϰR������Uoq�9�Bz��V��)N4��i�R���M���_3%-��ԃ�܆���)[����܁�Ն>s��Tj-�c@��8|�ZRߙ��Q��jC���Ką����_��?�3�緎di.���-f�}� ���щ�v��W����.��EXH<{mm�ľ#G�'N�,��7� �py�{�m����������5����(���NK�l]��QY˞�	���s���Cƣ��_�U7�k+��k�
ˇT����w�?b@�m����s�q~������� ����n�.сi�f@�囪����b��d�gH�=��������݅3���Ht�˼�0%�F�b.��cɿ�uz��S���zxh晡��|��yu)s
yC����#|T��}�.�U�?�]{A1�2Q-oV�>��ej��4�G+&�a�y�t�м�7jyh#*ea
p&���T\��vŝ�˗�_���o�w�B�E�(	iL�d <6^£��D�Ғ������k�B�y�vf4z?��䞭���� �ӿ�	cS�k��c���ܐ_�z��r�Q����@��Ȼ,�K�3��.*�Ř�L��}���;�wW�e������*9�UJI
T1y��b,%r�ٿ�P~�g�$��͆5��&�z��NoC"
�	W\]�JRǀ� �p��Ydc��@X�zP�غ@k�����o��n&�3�x�áD&j8Ra^)t~�or���"�^2V\�XS_��䭀�&�"�ٕ0�',������!\ �Ĩ�/��R2����<z2;M(�(��up�I\���o�����px�,��#ϒݳ�ҟ>���Z�(V�̓����-n��")v���m�H�#2
ҧ�x[444 s9Z��&�:��F�Ǎ1s>� ��PI�����p��}���5�H=�R�7�9�G>O�XJ�Q	��V�)pD`�,���wd|��mhh(y�=h�c[�-1J �F��175��o�K�؂z�3"��$Z�k�C9��{u���_��yA�SR���S~ ��f�G�=S�Й��9�X!P���>�Wc�5�ű��:��y��Q+K�:Dּ�u{�����u������?ʗ�a��'ӕ��~"�[��O�΄_�U��f�Q	l�Uԙ�����~!:����If&��!�rU���׏��r��<�-L�g-�UZ	����=������ϧ,t-�l~!!�&Jy�H_ޔ��g��Y4)���ߖȢ46&/+/�w����'��(�����E�z�}��0S�3w�[�o\ahl�=��|�fz���+�����lP)	֩��3�����FS�K�!!��fQw�ȷ��AD� P��������M�r�P!����跫�hD�{��O�BV'Z�b����M���_�ʱ^�$O�~�9�p��3��:�2d\�-!H�:�9�	����p��)L	y]�l	HN"C��*��Q��x����(�-�����P��S�,��SF�VÉv49R >0��	w'��m�ů���LS8� �7J��u@�L���ݼ��z��:*�qJ��=l2j�:����t1�?o��D�ā ��g/1 �#��@|���$Q_ȿ����@�WG�3�y9)�#����^\����e�����Pi������Ӭ�!tj<��~���Eѵ����M��f�~�8/���֬ˬ�H'���3���6��h�h7r�����g�`R',��Ck|�B�a/r �?ܐ�*^��a�9X�?��cO�BVͪo,�5�X�.����6CDW�f�W�18p{^w��2�RG��%�����+'	�E&��§�:QI���$^�W�*�Q����3U���f$�g��#�J�/���:R{���#�Y^�W���˱���iV1������	��U݈��ޖhhD�2��P�CGN<ĭi���F��j�v[�?L�V4����E�j�K����6] ��X`Nygs$P�6#n-��r��w��4k��c(��ܻ�h�m�D��>��5�U��Ӧ�6�e�~6�/�i�r�M�**1{��R��%3�90kA���ˬ���C�"e�v٠��qc�f��ؘ�#��W�Ǽ�Q���VqnY�O��\�vԺ���!��3BX�y����Ix�&�AT�.�kK�;;;,,*�t�p�R�Xxc��H�`<_������fJ�˜ aL̈́�J�fC���Ø�Г>~��Y�>���OB��b�o���\p�{�A���*2��A
����xl �q��1}���_ACd�SГ��\�(\�r�_�*� �s�G��rt K�^���_���K����!ņf���5�D�j"0Sv[m�".�>��#F׽rď	�2PY~�>S ��x!P�/��F�S� �A�Q6Z����J��������J�D;�� �������'$e�r͚�b��YoF-J�Nɤ�v���ј�^׹�J��F��������䷵���jp��=��.��XY$�"�]Ĭ�F���H@B�FH��Ӣ��)�ׯ�`Mr�����w���vn
 L �?Dl��I�3�&�F���Q9�0�����2/
~wɄ�U�*�#����wJk0�ۿ��ܜ�Wm0v~�2�`���j�O(UJ�����m'�`�p��#�u�"ȅ�-��io ���F����F��Ҋ���2���2�E�+��X_���]&kQ�^D�(���N��)	"��8�)P^71�Fh-��*�z9D<7n],
_�������x1��oe}�r��EO�)�d`��P3pQ�$��"�����g �}���B��BT_5������%�:&��������ќ�!V��{�K���F��Q�;j=e.��4MZ�
��G�~}b��u.��d�B	�^J�N���o�,@ܟ�e��X��4[���q=f)ҹ/ѐ �JՂ)+��H�����ˤʠ���HT���Z9H������D������hP¥W��z|&�S��fc��8����4�A���r�vb�����@����fس�6(��k+�ɒP����gH5]wD'�j�8�k��ü�';��EL��Tɚ��zb�[P�ʺ��l��{�^lN��E]�g�x*��CC���d�w���#�	%��_���X&��*��;�\�"D�,?�d��ѿ�ʧ uY��^(V~-?p�L� :�wǵ��t�/HFf���h�p��+�d@(!��]����L�����ǌ���O��A�܌��l`:�@���,?
�iVz���9��b���
��Bsj�mt缿uUl?%�h�z�����]��7"�碞��
���%���/�GJL�<��D0��$���b J	���G�(�62�Umn�%m5%p֎C�l 0�\[[�����),k����j�ݶ�)�&�?�A��ǅ��:k+jY&�ew�e�`�������D!��E.D5�P�<<�Ɯ&��y�j(��/%���������nQ�^Ψm8���C�L�
~
��a�u��s}�x%�E*�n�cS2|ٸ��G�[R���#��0D	�a`�`��d��4H�py^��5TF� �=� P���4#����Ğk� �y�	�{�̰���X:�Wg㉊���rm`�5m��S�+5��b[��i�A�|��k��%�:?��i�Aj�%�vd4����6+�2<k�0��W�F�7�z"6"�Z�C�-�����Ӭ��?�т·^�j~��y¾�����䇞�,y8ý������SGG1�~|$�i����ĉ�
�i�xM���Z�� T�n+..n�Q�v�;��UU�?�RT�0%*��ׇJ��=Q)P�ۥ)N�+^��hG܏k�L��0�Q�~�, ���#T?±��wM������:�~����"���	0�x�E�2�f����n��m��T2k��LC���&>m�>88��MK�D�楨�d��G�I��`ֆi�Z�[b9<8ݣ	�����,�AT��1���*a��
�6�O�3�Bxڔ���"Kf��]�!ԭ��5�����vy���)x�����s���Ƶ�w3=a��k�+���N���!�w!dd䉙��������zeA˟D�ա:C87� a]�Y+�59B�?'�SQ����ɼ����W�` �_T{�y�DK������\EzB�󥻞Q��S0�k�!�C.L|�%�K	T�$	:�9��S�����9"�Ƽ��i��L�����b��#$�:�s&@��E|�ɔ���yt��|ٷ��*����z�IS}G�'�Z���^4����l!��f	Ԇ8�����s�fQ�[w	�\+�^����3��s�3�&�o�B���n�N��B@���6�@_�p����I(Ds��F�wM �-�-d�ED�B��uo��ΖM�4L㍢�B�G������mGe�3�J�]0lW�#%r��M�ێ��=�����L��q�c�f�,M%��i�Q)3N�m�s):,Ǻ�[_��w�&?��%"��`��ZN�Uq�܌K ܪ���0LaQ��џ�u��P�K/������r�_ƴU��@���2����#�Y~Y
�o�E��aow�xW�ZTC�Fv=y��+5�b8����g%���RiP+�������_��z� �!�M�b��.�֔�x&�3A�	R^�����21��f��,�0��Ǻ��v�q���N�����]���H����?�,/"�0� ]ٲuW��]`O�
��`���֌}̱c�P|v��| _p�D�KB0[$�Ƈ6��g�~/�T�l���7�r������H�&_ַ�T{yո?oeU�a�y�6���0���8#7-�9�]j,��x��Zse��h�ќp�i��AU���:�X,����������/4�^���}�=ܨ���%T�C�u�4���=[v���u-�����C��̞��������А�N[��E�ק �U��\�5�&�h��+g`
i�z =~��j�f��j!����5VA*y�3/�::T����W����8�3��XI*�ZԢH!pZP�Q����,�h��p$ھ�Q��Z��:EDy(���lg��|�� '''���Z����~G��B盋xt�&.k5��w���SA��mZ1���t��N�x�?}�k9������CE�}��@�6R�,dԳ���Ϙw�=��k�ei�$���o_���厐L����~�N�����%%21^A��ݤ߇��
9���b��aᕠ���}ŇN?�8F�|�թ�q^�I�eO����
��H�LD��lֹ�8������D����͛���*���.�}�X���rk�	�ebWfE&���8��r$?K�*.}��o�l��al���%؏��Om
ND�(�L�����7MkX>@�4��_�AP%�˗B�l	�R��V���"�����-��H��G���riSr�V�>
w
�>��d����f��
ħ7'`3筡,A� ����J���CZ*iz�ݕ�[�r��޷ȇ=�M&�t20�PDv�|
h #�.�����ؤ��3X	�O�(�`=�I0jʬS���쌟X��XaC�JEAc&(�}���t���Ͼ���AW73����;��y8J���,Y���}$��v��x�d�W��N�U�0�q[��{��uS�֥sZ�
�>x�XGb�c]��&��b����n%�Y��A��Ƹ�R*� BI��/��=������P{V�w߶�%�Wu* b�j���4�������2��p�Key����I���%�U�p�5/���5e���<~U��m
�.�c�Ͼwص��A�e���Ä�,���Y�����Ě��w���3U�����*Q"n�˘�ꟗ�
3�d�09k��-�z������_��Ꝗ��¿�U�Kqw�KGE����']���{�<�y�a�'Y��	�O�?�eT�k�>�(X���2��(�-��-�-]Ʀ;�u��nAR�i�J��w���y�a�������;k�k��}�q^���-{=���iS&a��B����	<Q���7	�#S�b�o�����v,�L<����Z ����Q��?���>�5^ꠠ:�Kq�H YDh�9W��0���f٨ '�E_=���r������v��1,x{���/&��s&L�;�*�H_/I`��NŲ�y���ǻ������u*<��a��}><���yy�bb���r�_�62�{,&:RW�����؉�K�YjY�ϳ �
�ω�R��� �*�[_uEE�J�I�=�*�ޖ�(��:��>r:�qN�
��F���[�uF��͆���)`��0_����s������7<H&����Ǿ�u}�\��ŋVPc�۟�6o�h����y�-\�����޸�����?��������j����[7��o��STR��v�."!t48Ji�9��"Q�^)�Y��4Z�{_P�����FQH2���)op��l�}�C1�)�#c-������x<ĸ�B��oZXPth%��-\��=�sv
����-C<dw�E���ޞ�w|�����o
:����l���p������\�ZUll�fu�����o�MN�ǖF�'��� m����xw�^�k��\We.+���.)GURJ1Rg��pH�(�Kz~�X��az�͜+`�$++U�t�/ɑ�e�g_�ń9�.*�C�#4��A�t�ӏ%A��#q�^�n֩����xsrꑿ�]�U�������>�Q���;������J2����|5�p�V�52>��fO���f5�K*�����H1^�4*#�̜�L,:��6��p{e�Z�on�D���<�����&N�.}I�,������Ɔ�CuO��m�\?��u�����V
S
��CIד!�	W�_�ÿ��(6�¶vr��-�e����S��7t}e5�N��{��J��pk'�fF��FM�*�r��3	g��{9���:U�fȍ�i�Q��U9n��h�ʥ�^�u8V�iG�R��I��9;;��D�V����Y����-uz��6�]���3ڑDgg���v����Y�����=vA|��9��?]!�.r=��X���(���7�xFFn�Mz�y9˗�Qw69�
n�Nŷ�����헤���s�P!�&��=���7kw�n�t�G�n�������{��Ց���-,UmճN�kac�3[�5K{�[7�>�҈��F*G'D�D�cd��R��)��Z��=�vT���U����[_0�.Un��JN��@�1�k�7ӷzrp��hG#��Yzc�oBl��
��7�f��������[8�L�̭%�6��G�G�5�2����S�[�w���Ox�'�Pw�!a����'eͮ"-��z�������W^N�ξ�)c$
�n�*��dzA+}C����w�\�����P�G���{�j��-�'O��:N:�>~�w52��A!Np�|��R$���>�$9B��U�;g���;о��U�^7�:>�-_����F�V�U+$�}��p8�s�;I��7
n�wqt�H[$v�O��y�&ϐ��%|f������|���AC ��K��ѩ�������ڏ���-r��>т.>���G̸��5�w5�4����k5y5�%sg������n�x�5Ę�W����IP�Uu��R��L�T�q-�5�b�0��x�)PXW&�^�3x"�T����V�)OIY�d���D���#�	�6̦�_�E��=�=S"x����"=VlR5.�&�)x�G��V:5aU.��l�|��
E��{�U�r��~h!l�F]S3~ww������ё�c�Gg�!l�)���<��J�%SFM�l���s,��^-@�Z�%��p]E����CM���u�ց�,�jj�՜3�H梈�{R�
�KH��7�����F����Eb��M��X��K�/i*�Þ�R��Xb��O�: x��[K�����xOU�:�ZZǅ&G��$a��Q�'�,��а�P&$$����;����$���iak��mY����9�iY��d�T��OII	џK��Z4��KT��k� K�"�c$qW��N�|j�7�O�\�ҫ�9cbbr���� J..��;v6�_r�G��B��$$E#�qJ�,JE��Q�	�����ND#����+r?;�Of�WiO7x0h�Jǭ8lS����I~u�A�J�H��>uY�)�_��
���&�*b`U�Ɔմ��En^�pW�ҎȬ��^�����vi�'9���eH�$%Y9�!�}�]�Zr� �oR��75֪c�6�u�hG��k���.��)3�6��5�oº��_���i�IAKM]�}Y"㖢}WӬ|� �Q�0��k
?XW^qj��K4W�@�!~�_3��r�l*�aᛢG�RRRC�'{�::/[�Co"��!��_>:[r>҆�48�8�֍k�}���~�އ���W/U�}d`</2'&�8{�
��z'���0�����e���$Z��*��\�������2�*�������ݻ�i�߭A//M�{�daҖ��Շ��+��]���,b�xx������n	J�ɍ&q9��cn"�{uK&���ȳm��>;!ST���Y��jlll9`����}�t$bJ~�t��Ȉ��A���&0h�b�NSSS��$���TEY9������a�����>��L�D��9��_�K��U�K�7^��]p$ϒ3
���<c�yne��i���l�^}�+ҷ�+V��ܪe���S5l�V��H"���A�,Z>�!j�do69i锟mT5�����bJ��3	�T�+)Q��`ff
��QZZZ#��g<h�4TT�nnn	�n�&�)P��q+��Hd_��3>y򄕕��)�?m
e��.��@��pc����8W&�{�����~�n�3���6�訨��m�BB������+*T���jߝ��{5�_�ED|%d11�(7���(�S�}���;ݰ#4'+k%�om{[�ۻ	�e,I.��K�/���1��Jη��m����]�kz��k��#
��TGM{���D��6I�R򄭪�z܌�f��r�V�U�V�6?>�'�vW_{����<�j�99� xwN��'PPP  f8K^��$f���� /��gcg�5��H��jg��a����
˱�5G_#�k=Ë�{X��!tQ����pokad` a�P�T��2R,�| �� ;���84�p���O�pbif&���Y�~�����x�^�X�׀��L��䄖�VIL�� &�w�(�nh�b����pZWChy�n5P�j��پ�(&E�,D����e��j	�tɏ�`��5���)|�n���3�CCC�}$<P��ɟ����� v�\=�,;�O[��������ʊ��V:3s�A�������V& ��6ӹ7oc��t��KJJ��\+�w�W)\�7Q/ߒ���8o��
�q�Њ���m:�i2k��t_��gT6����&F���M!Hf���sК9�������	��`O�� o%9�P��� �o�����t��+������uβ�[.NWG��!���Hp�k2K�'����}ܰ�n%q��16��n���|H�BP�}_2O��W��'�H��u���
�p��k�d��}�l(��:rf��s�/����+��w憎?y<??�j>D.������f����%����.|s3fr�L�����i%{�R�������`�F�;m���E���*7�y�p4�&�H�3`YԐ	 ��bXJF���R��œt'S����]�,��x��o�<ݟsh��3Q�mR�   v	������Ϟ��	P��S6��N���S{�s����&�
��h����.[I0E�_�]Q��YާY�5:j�q:�7��NM�E b���,영J~BD427�EfX�'�%j���IY#�����gt��z ^��D�7w2x��D�;$w��OM�t�NM������n���ޔ��Q���}�v���G����?��Jg5^�����2�B�|Mz�GSs|}���J�%d��/^ǭ$b�5� �����c��l\DXy2�u�999R����l��쭝�^5����2�[����^6^�"ۂs����~�6��q'�����&G��.�D��\&0�2yJV�f5�F�9���V"�#�0���^�:��j�59�ӯ������ J���i�㱞����"K�u�״�4sOh;��	H���g�Ļ��h��y�3��f<�!U�aV�!
.S��р,��4��^�]���oR�����_;�n�����SPP �+j|2J��`~�lד;1�Yrk`�/�n�N��P�q�*羖%���Ex7̫{���9�? }�{�#��z#/-8�<�tM�;��E0/� 6=]�z�H�`ϱ���A�&D~��l������tfx��5;9M�8}L�[ �ZAY_�����0��l��O���Rlv��)�	,J�kq�����u�pN$Ѥ�p�·���j��7HUTUu�b��ʅ�(�?95F?n0� !�lhЭsٮ��q_�+�,����R� �x(Q	��B�n]�ˌ��єCLIիp/e�.��Y��bf]9D;0���a���J����'��Ў��<�l�$-�z���C8f��8�.z]��kC���y_8!�c��©���{�T^[�["�&��L���;÷����tT }hx8���PBf�E��%�)-��-�E0�
���gg��<��x�	'�W��w�Z����Y�l�a~z��	�����?��7z��7��ր�݉�}7���`T�vL��^������mc�ՠ՝��@�;'�dOB�
��ߩ���b���x�GJ
q2��(�6>����T���t��p#��	6`���t�n��)9bn�"}������cb�4l��t/K�������1`�H}���T~(Σ,��y���B����/�i��^�� R�	(�F�QWV6t�T�e��h��@�@] hece5뎦%�$���E��dm����Ш�� `h@�YBg����
P���1�N��z��ϑ���Ȭ+���������q{�6m�������MU0�aL��v�����ր�pXw^��9r��۵�W�X�^'�j�r��z��ު�ۓ#��\'��b��ml����M��>�*+?Ds	�|x��@���g�l����q��ۭ�-W���l,�����y�2�CPI��+����wV����F���r���N��x3�_+�CsX[֔<2Ask�
n!���rr8e^�u��J���]�s��#��̵��`f׵$�%�fj�&�$~�R�S�.�f �� 9?�v�ƕ��!JkS���oa�������������r#O�%^�
�����g�Q�1̝m23�3hZ�������%�`m4�ړ����f�Z�/땵[{����{�՛͊�J�(���*w�ޯr��ʃ��ݹr�������Y8����"��t���˽��@�iun]�P��<�+��$=^W���i�a�}�e�Zk���Ҩ��Si+rc�MStG��l�5���0�mJ�p���S�v�dh�#�(���%�س���GAn�\�wZe�v��2�L�����Z�j����ڽE����OT��2��h����o��3�nf�����c�>lc��׾���a�$P�~�1tJڄ`��_��_%hhh"��/�e�1z0��	c��KH�Mű��D���:F^*�����~$0_���>i-X��Q�����J˳ -LW���O(6�36���څE�*��6�Om�֤���ʲ�A�*ߗ��y��3�1T�#������V�CrG^��g	��0Ej��������$� ��ol����J"Pxyy�WRۆ}��{�-ضwc��ss��ÈU���;M���;M�_b� ��S����V���g�c�M�0�m�⿘,yr��L�_�ە�B��v�i}2���p9��(M��(�K%�r���t�2F�A�Ɠ�u�}s�/O»Թ��h����%*�<R�y�ց��a�~���h�	zlՈ���v��4�0��Rϳ�����Ȩ(��D�k��eĩD�qO��8�n��(�	��Ž?��-�����#/����t��S��_�ө�X�<=�p[� r��ڰ{8��~1��mn-i 1*m߶�� �Γ:�+ЍL���w��6o|�jE�6��3�+���,�BӦ����*�+=łe=���W�$E)�n�G<ˁ���x+qPP��?�W��%����E���������`�cu�9p�w�j^���E�Na�;O �	`�j8�SUS˅B�677{K�=� 9���Y����(�e�
?� ����Y� -({͊#�OF�(��m�錖�#!wOע�,���t��J���a޲��|_9�F-��e%7م_dᛁV�t�y9�a���`aaVOl�y�rCF���𚊻;༵����z���������ϑ��ʒO��������k���$����������3���V@��
�2T���@��W�s���:X���\���������^QK��j�pl�$��чO(��ʻ��.�w{&�v�RG�c�H�z�7y�R/g���"��aR��P>cЁ]�W?�:h�/P78�L�ꈋ�o��(7o8| �~n�}��e'g��=��Q=T,?a�8z�P��������uf׽���d����
�N|�xLCv����(������|ܹA&��^ȳ������>�I�i~C{�Q�w9�BEɹQ�!g(m���.��."q邩�<rc�.0�dk�0S	0$��"c�J������_9���,����K��c`����tRw긪��J	��7 ��]����؝�+���4�Íq\��ۨ7�ϴTT�#+���|y�2�4F�onڟ�Q!��{��{ɾk���U����"�4iqѨ@�A�j֫q ���57���Ӕ�~$�K��4Su���5$�̻�鞍W��?���L�asG��K�N{2O�΀��aJ�����?*�7��r�����`W��(ڽ��7$$�[^�x����f���Ɖ����@��o�Y�H�3�*/W�5�$Z#~d00:ʞ���i,�<O�`����
��-ۙz�~��&���e*���%�4�����AA�::���X>w��0����f*�Ę������P���Ǯӄ@K[)p�����e����PH�7"�8x/��UV�7F/���[��
3%�a�\��<+π���	@++�&\��KlN�;�b�BݬI� �225ͫ�愲|����Ƒ��^qG�\rn}}}����F]��}���Mk}�U�YX��Ǌ��OW�k�:�� ���8"q~H?_����T��� T6�]�F��D��p�vd�+��u>���|IU.ô��P�!��ڕX⳩��U��%,7r�;VH5l��X��G��u~�|ii	�v��z����:���5����8?#t�Gz/��i�:F�y5������{�Ą;�w]R�u�~${����������K|a�ė]��~Z���v�1`�lmG~s羃"d�d�i��z�]�	Q��c�P��P�u���j����򖱜����CX�0<�Y�u���4��2}�\��[u.%��� J�h�;f�ѳ����9sQC�z=�?v��b"����6+��#�.ųg�� [�s�����u�	��G�|j**�߄l\��V�H̼� It�~��y���'�'{?Ьs�G�aq��[��n���ɒ{���Eo���Aƃ=a�}�|�&q6����ç$Gz�1����������>�~�z���4hI�#�G���+C��>�Z�~�_y�땋�D��xs�R�q��2M׃��A�`��X�6�������
��|M�EM�0�¦]f=0�r>��(3�Թ�#X�:> �Ç��h�L����AS��=J"i��7�װsbڡ�Bҷ����N�g�'b�ė����5}d�i��KS#~$a,{���MtU��CM�0qOOO)9���Ł�p=���֩2&&��т���q�g�F]@��>��Ѐ�QT$o�p0Z܁���3�ey�l%4�u���4��b���ʨ���_,ܞt�!�7^�R�~9�X�h�������>~���h�ѫ���K�0
4���c�>� ����pJ�Dv�!�� ����OZ�¼IkK�ul���~�!����y�\糢����-xS��#/�ꡗ����NWӘ1��"U�L�b�z ���"��\�}_��\�tG����ԥ*`v������n_����`�Q�x����iqG��`�UD�T
����zV&�gsLѾ�l��ΛZ��M��_�<�?<t���\,s4����n܍7m���	U��)D����	K�T|�����8�]M-����!O>��ob���l����`2���v;��	�<��`�/	ũ�����x��i��ٹB��92eۉ }Pl�[D��U�z�(�䭌�#��]kDg��*��K� ���)|���D��,����om���; ��������n~X���?�X@7;�=^�4C2�5Q��x��l�@��i���e���eT��L���3�:�w�E������w�oqT?{�v���kӴ�ZQ�.+��F�թH����zu���oʊ�2�z ���1K�Ôz6���Jh�J%(,l����a�c��������]T1��׍3���>J�j<����-08��3���>��F3���ޱ��ۣ�z���Υ�����.�O�A%����:6��6�X�J��'O��;���V����S+mg'&&pIʼ.ܧ�'����4����]/����Q¯3����L(��߷}�~0��.*��?L�ɫ���[��~�H�4�o­RoRn>�����(B�&d���cmqh�nb�@�Z�*��jy9�%%Ox�0 �#^"�r��o6��i��TW�����ڄ'3<�����;S3��;������s���t<���Q�]�k�^��?4&�deNI�][�K�F�0�]	�4�߇Zmz�18.O-����@��M"W��fs��v���陇��U�4,���sKZ!��1Z�j�$hj ����z���M��!��җ<p6-33�i���^!U�;�v��Ϩ���c=��~�6�9h��̷gO�sT'����;�WD�2R�t&Ij�vȺHD��	s+x�ކ�����rTh'a���?�C����Fkc��U�`r��(�5��S.lT_UO����)pQ;��+���LߌW�CC��z(�&���7GKK���l����}P������D�$X��O��}�4�����u^vQ�mY� ���xu��C:�#�l'uTJ��%��0ڟ�y�uE�h���`���G�g���'#4���银��˞���`_Ԉ��ح'�A��g�S6.��3�N���v���w:*엺×P���Gi((D�#�o���QW�Cp�Lۀ�A�OMOOs�����/��LT��1�{;���ZY�� �ڟ����Tu��b�,���Q&^�-�E�T��խ5�;odSx5�� ��� �X�g��&3�����P�i$��y�4Yp���՚�Ml�?���h���'T$nI{Q9�Ϙ|��¥�oZrz��s�W�ֿ��I��ߓ�:��&7}����95ŷ�BM�*Z�O�"�<8(��=;�C�����`�&������q�������-�p�U�����Ca+#�!���T5���-{餦^;��(��C��uU��� ��z���*`)cI��-	��P�^��3��9W��i[h6_��;£xSG���%"�N;�����hk�^O>X0��V���l�u��5LP�Lی������z�Q�ާ�.���_~$jvvv+S����#���C�v�fΈ�����<C�2}х+ � �s��N.����YS��g��:�ji n���IHZ���2���S���[��Z'�:�ZZZ��s����[��l�e��jnn5�/5����B�^Yuuu�5���O4xT�q=���`a~��uj�~?m�f��]	>�kk�~�?�:�l�����G�e"�|/x�-��p�\+�ADT�勁�+6���:������g��ԁM�==���4��k��


v�.8xgM�O���@<4a�G���!J�Ǹ����J m�����Yb���ȯXCl�/IɀG�:�K=q/ `tl5���"��jѵ�ߚG1Ϛʂ��Jػ�56EC1��~4S�:�B�7����Ƀ���	%�H����Q�!(wg�����\���eea�1/@_KIF�n�kk'rss/rrR�.����9��cS��*�$�����N�� �g���<��	��0����^�XXݛ�=k�^����RvwwY�v� �����K;h@:���P�����Z/ ;�2w���gsI���T,Z�/�^sD�Of���Y���0G|�v����W���}��v6�N��&I���VF��o߄��>�p]/S6}�/ɦ�f+������"J5O��z{���ݣ���<���h���j���Â��]]�����d�=:�x��-��������{>�#S룠�R�b�{��X6�>��y �N��
�����c*���r�ʔ==�����9<�����9	�����畇|������p�P����Im�Q`0i���׹^C�Uae2o�&(���?(����g������$P��6!�(73X�镁���.b�a`}��6Y�|����-A�n<�����:�"J����53�f8� N��b2@A���LMΠ��'v��\�-7��4�o��Mk.���>����y2��q�E���q"]��K'1�Oξq/��<=�1E�v�s,맿�)��sea��>���v��ڛE�+�������
�hF@&8�}�7'c8��v��J��Z���{�1@���
t�Ʌ�j�э�h�����@ tU���;��Ʃ��Rn��G<����'�f��M�mQB�,b=(C�V�	ڸ����{`���fa��Haͧ�6����é�O�ǃ��7%�8V��+W����1%jsue^��$��O�	C��3���嫴*�3�d��c*����[?Z�g
j��V\��ח(wbei���"�(�2P��0PW�IT���w�T��YdD4,GXwc	;^{���.�+&�4{V�C#i��K
L�k���ְ��?Ty�um70��j�k@M�y�<ESC6�I�I����їm��ꨡ�P�b����I�bnt��^�/��!w��坓�M�����tgY�k�M�*�|��p�����p�j�����뀭�M)+)凢jt?�������ʿb���[���g�ї]y���(�_1<��� F��q8����g��Gf�����+��ޮ�~�;�u,�h&�h{f,��#�,���vh� ��N��g3PW��W:�
��pV�Lk��\�:5�Ž%��=�7XW���:�)�r0����n�T~���*����U����+/�{{ӻ���q��,���c��#e�u�Pm�������2�}4�~�~c#{�§����j7|e�*؋B�o��!�ѽ��}gμ��w9�.��ҚӍ��?oݱ��?<�^?Ђ�備�Ú1�'�5���5����NqG�e.��ۛy�ô���Foc	k����w>�>*:tT�A^�����V�W[n֗'r���4w�xoV �^]J
HD���0ʛ�1p¸�Cg�p~��u��-vVQ�USK^�l�z@��]�`����!¹��*�NJ�����F+����ᣠH��P���ѿR��^K�<��8�kB�s�cb�ĨX~Bme��Y�?V����z�c|�uR�������h��|���	��m�doL
�2I.��4���ݛ���CCC?� L9,���w�:�	����:#����n��J��l�X*�՛�$���A;L�� �?����g��a
;]BN�]1��J�q�:�K�����Le�-|֤J�{�_�l3a��?xܪp���6�~`����� p����=�4l����h�I�������ef�\c���|�de�D� %t�����=�s�F�k�}J�J�� ?ԡ�c��O�}&�4Q�
+�q�r���ćZ��@�^S}&, IʌKF����������������>�:'5�j֕Xȳ�j��H�/�)>^�peE�W� vY�r��$'^��S��U��s��rj����Q�{��E��=ٺ�J�B�V�ܧ ׃F�a'������9I�#F{��s�F���{���bB�i��gY��-,R<_��������eȳ ���aÄ�FR�K��g�E	%�ơ�BMZ��*��@�j��&g@SA����ZO��@��歮��]�#�f��/���E',�|��%e\����QN�g�x��KS}��1����T�.�a�1=����kpZk��~�+�F�gҜ�$�b����:R�x��V8��t�f�|�W��m�/Vu�1I2��vC�1��P9+L�+���3��d��D���Ţ�.�\�!��ii��=�Z�z����31<�0��E��T���)�?m�W���T�tKb�;�H�w8A���Eg�l�8S�i�L���z���ޚ�y�e�>�<C����1k�r ��a����@���:�. �p��J.l��f�rS��`S���><������n6QwZ���S|�Ol�t�G���#���3�Y0\��Vj��� �_��?���g�Q���eR�6���������AA�{�;Jm���ׯ��3M@<�C���Q
�
��5����ٯ�||�u
�ߥ�J��e��������>W=3��cNqG߼CM�")�c�4SV�vpxJX8Y��}
�Ĩ����ک��y��]�z6_���}X1�>�iD�5ǹ��k��r{<2�(��`�K�V~��w�oJFg�M��IZ	�V�c3� �U>��b�J�s�d�B�{-F�w�9mt�Z��?\�����?�������U��a�K�"�踧�'Ej��Z��v>=TG�����0���Ti�6��)��	�&R�S��V�����91B�E��Rr�{0[���}�� ��_�������x���4d��Wa��������:�qU���^���z�i'�>N��~�"�Y7�!��Roj'������}���닙����Q�W�c��JEb!�3FYC�>pz�~�t�����2���	Nڪ��_�u������N|s��))�\3,.$�:�Ų\`PfXł�����P��������h���8h?>�[��P�����8� g��r�t��Dy��&�Pqӿ�˳�,����;�+���R��R����8o� gj�P���Nu�N�p��I��G�'n��p6K�͐mޝ7��v���=���!q��h'v��v.˖���/ٱ�"ۻs��X��[&��(�F�{/L{�\R�x|��( T�tvG��g)���V��}>�W���E۾�D��.B%%��$.��w^����������>������CEțC3�Zt�c&~�Cs&���t��y�����#rH��R��܀C	l�4p+b>F�F�&hk�ϒx3����9��\�V��}�Ք	����4����K'R�Bv�fv@�T'.�����T�q������8=�!���s��ٯ�7����]�5���""x��_e\�+W됷i|>S��bqi���OȒ��F���I�|[T��'���>�����i�
�'����~���*PW =�?�al�.o[�,G	��D�+Ue�'��K=i��$~ەL[h	�磏�z�F�ISe��=���õ��^~6��.�Jˍ
e��[Y����)b'�wnr1jf-˭xȈ����JG�)�u�7���C����bᕤG����ߩ�85��} `*I�|��z�J!7�={��Pa�$�
���2KC����4#4�X�-uowA`�$��m|*=�7�Bn��v#E�A�ctp2 jژ��M���[ �*����'�1�Q�"�R�!�)9u٘�f+�@R�y���6�ރ1�� 9�d� �l���wnzڀdW�qGUa�Q2�,yM�@��P��|a�]���B�3�p�N]��@a�!!i�Jܣk�����T����\�y_Q���H�k�a���N۫���pߛ��}�+�aA���Ba���b�;{C�=;(�ET�W��qq�<� J��6+^=��x޸?���$}PR����R�ˬ���E۵
{t�Mz�:KV��!$��(�
�f\��֐.;?��<~��Q���]��^{H[�5��*���u[$0���|���Kvo���|�*��^�g<�x����=�~2lq�d:@�5�
2���K�Th/׬��\)�&!Ù�i9��G�R��w	����='O"�(��m�9�C�"���>�0�x/s��#�O�[,���{.�)0�Bя�c�W���^3��q/�m
����<h�S*HZ��p�R�QǠ�`3����"�^���X��5} �u�n�	��D�>� �q���GY�s�S��X_F%FIq?�Ow?�I�p �ͥ��N�b\#h��{ڏ��geM?��5��3:�-K��q��K\2�IͲ�p��&?C���\�&�!E�o$�^�%ց6�R����4��8XE���:���Jۖ(;6"`��l��)���pA���e���o��u���Zn����[�$M�Z��X��Hr�kR��=&��56������=+2�;�K@��5>]0��s�
�R����X�JHZǵ�@��XN�� }T��+���S�[,�Zi�#昭.#HzM)�C���"�	�5�3T��L&��ĵc>^R|Uٚ���3�!�U�G�P�ּ��ACdp��� ",�a��/:��2�!_;�9LRk��(�)'�m�Y����=nڮӑ������>���h1�8�p'8c5T�=��k`Z��F��!�t����ՄmS�hR&�R�m���U��P#��S�i��<��m}`Yn�����k;�����=�����=%佗E_�ӻ�_��{w�}}R�����j�R�YV0hɪk�!A����^�iQ���Bz�QI��Ӛ�R�:��'���V�Ї����fش����-6��� i�|��A�K�Lę������hsq�WR�e;�����W�-��<��C�S����^R!��ِ�!	��醌(? �Ɏ�l�O�|��-��_� ���g�V/��zܔFg�f��xyB7����A-�h����\�TS'����<&�@]5�1�o��~5Xm��H��F�)�1�r=�P@=���@Kݔ�θ�L&���E#ōv��gwi:Y�5[E3���JO����l{�!\�׹��T�_��Rǐ��6+L5�h�A���v��!]r���>׭h
o�3���GQz�9�q�5��!B{k���Pg�br�h�v�5���93B�1Q�*uS��O��4ٓ���C���2�&�@P�yT�"�I�i"��"��]�kjڄ]Cm=�Ȼ�kw0;ʎ������Qɡ�v-|��~����nj�Wi�؅�����k>=���0x�ye7�E��p�����������:��ۅ�I�$��{܏�
QoǍΝ�OCiĐ9{Fj�dv��r��X��<Sc�����6L�w^�����(������_�����k�\>dx�pH�����Q�N!�f��1ރ��K0���`o�D��$���Jޢs��i�|;b��r�oDPV�+�y�o�.8â�W�L8�JY[ȁz������>���OlxX�u�ɚWu���ܨ7;��}�Go��
$G<�����&R���������<i_r���	*��_�s�)D:F멿=��ޜ��Q�d�,���Y���\���hͅ`�~��P��W?ܷ�҆�ٮ$P;���0پ��q�	��n��B\允/���ՑdgP��S�RS����+�ӡ�PvQ
�p���X>���Zc���_j���U������E�+�E6yn95IQ��K�b��8M��i�d�K�Y��JA��U(�ڕT4�g�cB��OWj1[7z߱"La�4��mf�R܏����F��R�H���={��t����:4�jalj~wR�--U�J��%�!�R��Oź_]��߳�⣝�;h%����f�԰>�[��IP��R�S���+�A���d����
�~ ����aeg�m�mxv)\����xsT��먑^`F��O�$8���|�� �����X�wo��}�~ox����
m���=}����[Qy�D�ۥ\`&�s�����62��2E�9���5k[��.������n��p�� Wm�$~gW��W�'5��Dp?��g���<dP�5��_;dL�=Lo&��ٝa2����+^4�0��9D
"\�4�k�,�UحB�}{��i�GeBo�.�N�P�ᥑ�9�5R�,�?ڝ�/�c󍭕z\|%c���/_q/��Z��\r՛����~���^�����w�u�Q�E�����g�-A�>ri*gj�p�1�mZ���`�$��V~����˃;�A��7�5������y�����65�w�������W�G_r��Q`�F�IG8�6�b�\��o'��ɼ���O>�79DQ�ʗ7С����BЙ��\��?����eu>f�Ο~�����	+:�r�/�i}�ظ���򄓿�V��6=��^o�._:��>��|�ӳ6���q��ۢ��r�z%C�n{+ r�
��ӝ��|�9��8{���-C�"�uۓ�o������3���8�)O[EEzP�MY�V���|=�g���l��uH���Єߛ	��Ԡ��50�؟)1%�����(�~yARu��^)��n���_QX�y�aN����$.�ͬ��O�,����6�>O�����Ln�j�]"#����Q���t�5d��;s~��e���Gg��������dy�u�a���P�,-9h�F�7E��m�����.W�G%��ްb@ƨ�;��F�컗b#x��K���^�J����*>hX�^��sfMo�,��"��x�Cb�`�u�8&����5��`�m�^��Z�Չ�L��.�8�>{��q�A���{!�q� 'pw�M��f�雝�S��[����Ce�[^��O�DAS�Mo�:[z�V��M��>V��Ql�I쇰#Ѩ\���K�ښĢn5���G�g��A7C:�.�"\�<<y�6�u��uD���G��2Y��ʐ�*[�yk �A�#lw��a�˜^P
D��`��`��?&�:,��{�%TJE@Z@D��	�	A�!�F�������������w��C��ҙ�<{����ko�[�7br+ѕK�I��%~�9���7{����t2��M���j�ь��s���Ga��5�a���y
�����-�m4	C��[�^=�:�i��5�����H����Y1Z|���$o�� yJ���R��I���Qy'%�
Do�D�/ ~� 6�8Lf&�?ntlb:�z�W�jX�����^R�`��F�~r!A �P⹹�Օ9�}d0q&���JH�.2m3���Vvܼ�1s$Ӡ���oJ9��*a�k�K#=�#2��&S����(���N�	�4�$FPEf)U�ޯ��}�Yr{�Ex�Q�K#�|�:���� �˿��ݝ�o���f��� J"3���k-��"�ۻE�0����4
��J6]��x}�~��v{���҉�M���xҫ@��-Y���͔�ez+��p 5���yr�v�/B�z?Ed9�2�]�ۙf5��T�@����2ԃk��Yӓ��c�	��S�"�"0Mn����>�.Z����:h�|Zé�+M�u�����;^��D�{�R1[]���y�{T��i��nY5�<j��t!�܉�:=�����k��9L��*fʽ?Xk��cq3	]~J��by�d�^v��|r��&��<pSPa���/Q>kn?�iz!�����U��M�u&j���ub��@����B=:���p�|�{�a�$��t/��x���j)~q�j�\]��i�m�5O��L�M�*���jq�1��	?BqMN,�g����d��_��v�kqd�aZ#<��̭�#�`�y3-^�	2�B�OnQ�Zr�|q�p�,��i�I�C"�>&*�M����Siv�=(�$�~-k�X���CD�rU���/V18~<!/z#R�ҏ�ŰYQd�x@�ͬ�F�{��V4}0O��uXk'&c��V�9��B��N�^~��m���+�Gc��Vj%ϻ��dXi���E��Ztr��t<J�w����t]���\��	T&yr��ωA��7�Й�p6���A J`z�-���_�u��ݮN/����}�Q����j~3@?���FG�P�>bLm=_�)
��/��π��!��a�u3H˞�0 �iF&�����5�I���F��T��Zo,ܛ��Bt#5��sv̲ �&:�;�?͜<O�l��a�rԵ-#Y42J��V'�w/c�>� D/�:mŐƭ�X��$z�t��ޛ����JC������}��T�@�'4j:*��z�+(�Q�&��i���<�����zB�v\�_����dPVǭE��`}�%@j�b�]�4�T�{}\G'X�C��,$]��e��vJ�$���5�0��TT�0�8�O f{�e}5U�h��]�4���"��;8���un��9?����3�1���B:��m�>��HS�1*)Q�+�m�(J��[fz�Ұ�����4�~^{��-i��	_�_L��%0��A����d��O����������<�q����U�c�8��{y���"�	��s�nɂ�Sr��%��te�ի��&zUz�g\�'�uU�1dM�6��jON�-)dFf���W-�5P��}�lu��>P�kry'�hf1O7s@'���d#Һ%/��cN_��01�F*5��\'�+ǍU8^S�F?#.����.����ŔF4מh�"����H �P�I�H�4e�U יd:"��u��P�),�>%'7b�h>���������{7����E�����#��e-pa���C��0WfS5�3�!(��35k昈脁�{��P�t�F��ǔ_�"�X4�&h<e�l�"cV�k�.K���|A��������!�B{0�c�̨������UE��8~8���U��.�VO�ީ�14N�� Gr���?�&��;_ǹv}*�ޏ?������]���0���d�V#ze2���ǧ݌�	�����1�fk�l%U�K��~1=����9k� �36�ܚ>j�a��L����U��o��g�*;ײ@C3��#6s��^*�v�կn��uuؠ�>�Cj �$�A�i�pYe����a�����Z'OV� �ڗ�w��y�H�[�,�r~嘐ZO&M;J��⩆����w� ,�S���O��2Y[��A�번�~���E[�a����[��������qX���Wڃ[뺄���P��#,qg�A��h�i��J�<���M))KĠ��I>@�S�#�M)�tvOo��v;�n/y���\��9�P�u#in�ӗ�eW���-S��x��i��Q������I@=���١�����"[n���H�~���6m��An/��҅�')[�KV�u�Dzq��0�)7�W܆o�DP�����rz]��Z���n�$Gv�n9���d̂ >K���	�q9#{j�⹌��U\_z�=�K������B�
���l+�!-��bZx���Aj�11�����p�D%|�q0օ�}�v1Fb�q�5�MW��"��aL��N��h$<��A�>I���4u8:d��R�� ��QD䊧{��4,r�L�'2,P��9��xW����ʚ$r?u\�vs5A_,{b&]�V�l#��:��N>��|S#��e�i0U�ǉ�"A� �.]�ybf�l.CҧL�GD#��n��j��6��s^�/RUm��X��ɯĒ����&|�8ؔ; &]�]���N~P�c�x���Hc9���Ѵx��m���Sm�L��zm�Ǧ�=� p��.�)�[3���Z^X&r'����'��2�޴�/^�l��F5��ki�Ŷ�ӧ��n��E衯r���n^�����gզ���R�<a�#��u9��,���D1U�����iN�s b8��P�P!嶺7@!W�ɃϢ�K()��)w�ޚ��+5��(��χ6�(j�(H�4��O���=�B��*tWˬؕ��C�ΙF�D%S��u�OR����˚���IЫ�	��:$@}�0@r�<�F�c���᭳̔��u��ʻ��p%p��eA�}�.s����xjt{�c����>q�{>�/E�hA~y��ȗ��x�!�''+�l���w�������>�sؾ�����N^2J�7�Caä]
"�"�-J��b�WD=U�2OgT|w���d�������֏�u��nfy��C���P��L������TRV.�եA�^�W�&�!+�^M����/�Ψ�S��uM`i�ko'��?�O�fx$t�Ir���]����b��b\����J���s���R�|�P��rÿ����(˂�L;=Wq��7�D(����iOEg��>G�8��~��(�0����:P��z������ՖR#�7N��� �j��?���-�-i����E^P���vŐHx�VVK �ӏ���)}0�i=zE�s^/��Q>����׮��������G'�L�O*��;�2/-�*E�
�E�z�L1Y����W�-SV�]����)j�#}_Í����g���
����S�ٗ]���
Ր��By�÷���E6�����j�V>�4!����%����'�=��*�_P�����ӕ��۲RM�N�6G� ��
X� �ʳ�?x�4w���u4y s��d���zD�H_h2�o|�g��F������ŧ_�E?	5��0u+$:y�tU�cna��xm��a?du@"l�XL ������V�:��I�JOcC;�V���<�V�|N��{���`pjr���<9J3%|�E��ln�,.����bA}���D���v��>��#R�.���v5ݛ2 $�3
=͋�Z�M��kEN�xƁ��K��G��,9�C�+�:ɖRaĽW`�_˄�鹁m�ݻ�����ĴH`��� n�ɣDvFO�)-���è�ݸ>M��=�A.��~2��a�g-�FA�w޲�I�2���P� qyx�j�d�#��4�����]F��Fs�x�"ۥx�[��on'na��6 ��ppÏ�(��j���]�E�l���-�e��$
7l�Г�-��{����h�I����xZ�x]���rR=��#��WxȾ/^#4�h��Љ�#�,�O�<����"]�|��ջ����0p�n�atG������'Ϩ��`I;a�ٴ�R��,ٽ;=����:�Cn�J�(L�D��Xb=\<��=�N��@$
��H���N�}SͿ���e�&f��&�N�>�յ2�
'dkB1�������ov���O��ο݆WpU6�ַ6��Ano�d����t��͂�v������D+�Z���(IA�ĹC|�kTmgg���h���h�L�}w�y(4\pwd����F�*"8�>w�_��Źb�k��2P��b�vz�W�֎�PL����[��R�}��
_�aim�[� ��j묟]�V����nC�.�}�o#�f��AzZ�;���Q��t&������9L��e#M8ۮ�)��o����Ga#ѻ�Vw�q��������Jw@,�9��ҁw��q�'z,Z��D.�/�I`dO��~㩶wIskQP�!�)&�h�+�0y�}a(�"R����72��`�pP����H#DykdoHM:��w|�zA����x�y��Z/�
���r�͈���iR���eY��9`_پ��:��L���b����_p?:�k��u��� ]���d�&�ҫIt�2=dT�@~t�h��C��b��	e�^�D���h�$��o͑ԵF��{2#J�<xt�n"�H��J�ǿ��>��3�O�$(�-?E�U�A��).6�2�Zwk{N�W�d���m���b�N���"��&q�iw1MU�2�_i�8��_����dP0���bl��k�Z܌�~�s]��]t�	)���|!Uw�R�Cg~� �9�D�~;��@��c1=u*�o� ���Wa��ߨc�QGamW���D�o��¼��e���|��6������i+;"�_�s��DI.�������CbW|^�#-�Vt�o����
����(5���)Ga�sN�WJ�>q������8�ae�܋\8lT�?��L�䨕�������
�!�ш�&'�I�O����c,��[ S [��2�q�Ipq�q�j$8�EG��З}�_�}�I��L4���->m$D{k�T�������u"p��w�	]�/����G��T⊁��BM��H�Ν�_mÁ�:�{N���$_�Ȁ?oɗ��hZ�%�'�����M;��{/c��ˣ���Y�]���*��
O#1{�E���{t�`.�~��t�ݼl�)�k��٨'��ٞ7�C����%=	��q�V_ߓ���rB�Њ�F@6}�&���,�����[鋜��V6G���W�R����b%w{�%_�O�m ��Ԃ܁6�{:KC�h?�Um$\��_�����Fl.�+߽�����nƺ�A{{��p;}�J�3������L4�9 �Q�U�s�ԓ��]�"1Ҕ�����ޞ�ֳt���̚����ӱs�����nXC˛z��H��{{d@���DD"֖"e'�l�Tb}�8W=�P�ѽ����suC���DW&3��'|��LJ��fΓ3m���/�AԽ��LV��IFB#���6=M�cM��۱�V��ѡ.K���6|��  n�����{���x���Nh�z�o�j����� 6А��Av�b��ɺ����\��q~5��}�\�i�2��~h��$o�J�E��8��m�b��2c0c``�iD�����e���eϣn�#�e�+�4��k7�UQ�awI9�K	�w�f�dVw��]�����r�Ų�����ǝ'-�\i�v��đ�����ؽ�ir��E!��V�ȳ��Oe�r��!o�����?.{b9��	%�i���&l�z(��V	(S��@_�d:`�gb����>n
9<4yv�\�hf,|0����f+R �u�W��S�P=�+�i�4�|���=7_u�����梭��E��#���-u��F� BɞL��r]N�����&:/�eH�4HB�1y�p��|�E���p����~d�����*�yBehA�*��]�u0�X[n[;?��G'tl�M�s��}v��/,7�����+[�x��$o5
��p[�+��#���'�p[f�׏d~�M�o�bš�'$i	���]�m���rV�P��i�m7�� |b�F�
����ȼU>s5-ՐB����A޴ar� �LI��eՐ��Pc�vx�䄄��aw�8y���xӁ��1l>/v��Z���k�<i�e%�׌k���K�3*݌�ݻ�Tŧ�^D����%����ym�=�흸�����&v�ĕȽ�%%��O�\�	Q���Fd�I~�d�Faf�]�Ǖ��o�	�uăE8QK
+|�<R))�����K/�'�jOA�y�ec�?#�Dm�t'��C�o�a[1�]�z�	mפ���iRd�|���^G�>���j�آL
�d��=��o��	�GL��&l��\Z4k��cm���;J�������U��k�����'�������Ó��Y߯7+u���y$ʞP��'���R
�)�������G�I%�R2O��*E�84��q���j0d���s,!EJ�{G�k>�!>��'������`$��|�Ω�갭��^ciЌ�v�З�ѳKMs����\!�;�9
����Mr�9݉�?*��$O����C�����x�8�*$s��7��)�R�WOj4��|,�<#���l�D��7���#����;��D�*�ĩn߹4t��w"���_�;���s��A� b�fm�n�oq[v8��� ���\�%;�>՚�}X��t�+��8��:u��\Fg!��>0�.�=q*|���O.�x�����
���U���2�my�]Oy��8<Ulлxp�8�K3MUm3^��� ���"i��Q�L�[Ɵ��h���t�� x=4F�z�����ߧ�	E�m
f��޷����-D8̿H;�2�K�����QjNm��?��W�S�x��#�/Z����mҡɕ��Ϧ������Rcq��NH�՗6?��ǲ��x���p5��?�"/a�c)s?�����Q�_�<��j��ڝ\7��C�vު���R|6!��X�^g���&��[Ĵ;9P���0\��_��q��>�V���Wt�j�����w}�S�?����D�Nq�t^�L]�tÈ���cS��5�W���T8�/��}���N��ɝ�L������_�M�@8#:w��a���w�G���>W-�[�@��{a�%�౓E����ꔷ�dR2�T���ُ������*E&4F�n-o!�R��$?/@鞳ggL=�h������o�7�'�*����ר���c���ՔW�e��{D"��qc^`���$�ɸ����χ��������\��5Ѵ����������:����8Nw����t���,�'���("��Ę����_�Ta��r�S�V�\�1�w
h��7�G4��YG>9T�Xb�_�T
��æ5m����B�Z[���1��-����W�Ry���'�	�Q���6j i�3ٯ=���՚b}��;(+(ۓ�E]g��ކTI���=���$bnM]ǅ(<���&��0�/)��Sx;Ч�f���Թ�#>�B�hY�F˰�Ɠ� @.���UL[i7h[	�9&���4z�?����b�\.��o;��?Y����oL�sAن��[#�AEI[��
=&ZC�'~Y�۳��-s
�57y�+��!O{�ˬ��¿+ O��(0�	k�s�q�r�f?��55�md?Kn����׺rB٤�j�7������,��i U�W��)�=�u��U=�������f�h��v��q�JɩQ8-��S"�@n��UB��荅Ȼ0�l��"o}۽����i��o�����}c�l�M�W��f⠴�Kr�<t�a��b���$-m�8����38J��?S2�+i�?N^�Kx���m�Kl��a(����Z�0mIS������Ǘ����^m��u��.t��E�]>sU0FK�|���I�$6�\��F�**�E��:��ICp�u�
��\.%K7S�6�C�ԝs=�uX\���͆y�	���u��m�XZ�ȹ��&8_�0�:�0<2��c��4��fb�sb0��;������y������t��@����ĉ'��\hA�v0�S%__	��4�&Z�T���G�T�h�9bi�R�EkL�7�f�tkw��� �|%e`tOtj�v�3.��,Z���<p�zw�
x�B�VIi�����u��*1A+��0���,z9;e١Dє{3P(]�9���#`ҝ�W9�7�i�c&��@�vҾu��+~��寮o�c`GP�|���踢������/Yhj�>O��/�b�> Dv2��_y���2ҍK��d�������$���/��"ަO:P;�c��*�hEJ�dV�2oۖ���Ƒ�8Z��Kcg^r`$V_�w*�g��[�-�o#Jg��&�+�]�m�Y[��K��o[���F����+֑�.��ZU��%W3NR�SX�15��Z�Y�+������"L��j��'�9��&��n\F�"��mD�!�n/��N����)�F�����C��4��9:1�B�w���(6�o�tL0����e&]����3=ч�`O䙛��� ���t/�w,����S��M<�@O�p~�ύ�5�8�0_�f'��ё1hb�.�2����褘�r���#�5�ش��N	w�I˗����>��~*�Vt���O�t�)��m��`�`�\���!�
�]�,\���.7K��9�O�=ܕ61zv2�i��ΩYs~�^�<�������C=��+,.�M|*)S�/Gs�q*z�4c���
�سق쁠�OzͰ�eEn,�mR�� .����XbEr�J�+���Ku5�뛡�� q��f3.���E|	�k�X'�q<�vbz2_��CN��J+rDO��ػl�п{I��8��"����Г�rz�$�3n���s��A9�i���k�H��qGf�w��e�s,;��_.�b6�Oh�&兖���(� ��/�	G+d}�1"��]z����#���K�ȏ����3����\L}� �*�b�����o�I��\��ќ�	�K��K��߶N���,��H�vWn�f?��h<td�Y��<5�q�p�r�ݮ�W��3�љ\�:M�r��:϶�d�R=A�?Za,A�PR��bcx,pl��64 	͚c����Fh2_�kn�f�λ>=8�B��p�����`nÌ�}��F	��Y7�����c�w�n"�an 3�׽��'1��R��OKj����Gj=^�qs�����]a��{�¯��ZZ�;QK��#RUƄ�GU�A$���4�� bxY<�\��wю��ej�6�t
����%���MW$�[�����"�'|OBa¾�3ޘ\���#�ۆ^����4##!4ك�
�}*�ɻ��-�z�o;�(ho�:˨�#�sM{`d��c�h���j) ��߸�uYؤ\.i.���D���'.��'2^~@�6� (�($!��7*u�:��f�.�k����Q��"��e�l���p����!0��^��jn-�e
��50yv�c�d�F������g���5�5�E�\��X>���v����ȍd�'<ֲOR�:V�������V�50:�������$����@}l�C��ܚ3Z/��\���X���1�`���{'ю�/����ƖfF��lL>π�QO�̾ۙ��䨧�1޿/}��SŢ(x-�4��jy�bc�Z����?��IJ�>���A	�Ԋ�醑���䐞���l���Öƨ�Ƒ��,����^m6�"�ݾx M���������Q����B�&�g�[�J	5mc瑾2�Ɍ�<S�߭X��Gm���^����m�X����䑎��W�,~����p�G�
�S����wa����:L�N���B��U��s)����_L᭾=�T�j�"o�>Y�;umKe!t�-֌�;�[���
����$��MeˊLXM����鲑�h��`(�ZU��]�r�+D�0���K5	���"��UZD�)\E�E�V:����c�I����a#U٪'�P��������6E��g.�U��(�*�g�O-U���G��h��s �ψ�8�|J�H���t}0�f|��M������>�z���۸���q�,�m�E��H�|�|l��V\�� /�Cdy��k�j�J����C���ޖ���m�'�c�U� ���dÈŁ� l'7U��7���7�TL�#�$ܷ>��_��[��G���0-T&�-�D�w���顂���չ �N�4Q�@�s=���>�zp��"Z{�]4W����)G���cL�)��R>� �#dP�Ğ5Ĭu�Z�߈�X�@�c�����"��A7�E؞���ҳ SE�kw���Z����wf����|����r/����kI9B�	v��8]�N�\�ͳ��ֆ-��jMs���lK���W�E1�U��'B�\)�k�.��E��Ϩ�.ࢾ.���m�#eM"�\���83%�����,�f4�Ѡ�KI���l��.�|N�yQ�D=B���~��u�=xQu�� :�\+c����!Rj�V��Ϭ�h�-�&6�z�����'�	�!`v6V��;ݠ�?T�J���(\�]~P��`������&�ɯ�p��M3^��n{N^�Q
H�^96���7�2G����њ+)�!��餩.߫����\���=�P���C]���,2�P�=�8I&������3�iW0N��a��If��Y�F:@|Y$�cy��Q�ʭ+�퉻�ٛ|(�e��6��mQ�ewxI�ݮ��I�x�w�x��ncC���8�u�9���I1��`�~�8����a�2@�>W�N�K���Tl(�P2� �ġ�c��{5��K���O�w���WG(P��KM2���*J��7�������iF�D�ܡцe�Ă#�nF9/��߇\�����G��^���e��{�ts�|�[E���쎐*�tY�=S���h�2��8�Kx�n�G�؁]�7�;�E����ibq������6�0�* 2\{�q��Kx��pw��Gh����k'Nz���L9�NV�-�o�2�����=�J�,Т�a!�^�V��Jo�(��nmf�8�:�K�F�AA6�>г��Lg�����\�n���Z;�����G� ���j/G��@��];��S�[�;�ZJ�b1u��T2�[0%��A�?b���R�w��$�bNs�%A�r�l�l��&ERlk�z�:�'�G�)��6�OG��3�ׯ�>��H���(�aoKn�?�\ݰ�H��kl]<m�0X��v�ߊ�F�$��yW)�ę�k���[�
�3�1�&�@:$-	�]j<���=<�3[S��#��3I��"�b��׃�oxY�[�c.
���ҾG��wA��,V�*�g�Tv�:��M�S�?�K������#L����M�4��sݽ�cw�t�f���sd�tS"�w��#��ܼ����E��P�u^C	��6Iu�SUl�V�E����>�[�m	�������̏��M3\<�I�u��l���Uk���ͻ��Y��T|R��\~��jJ��� @��ģ���H(c�؄�~0��%�ڳ�n��~�t�+�Q��R�_BT�o?�G�C�+�>��q
'7b�-~��Z�x���l��Z2�*�g��(���ٕC)D�)Q���	���I������f�{�o�X[1��Ǳ� �q�~�*H��ud7�2|~�%H� @��4kr��ԅN�.��̹?���{���[.m,$N�+�a��6�n/ ����f]�;d�n���M��N�A ȝ�5���xW�.&Tv��	��.�B{�8�!d+S�[�\ V��
�c��8^9/�ڄB�oz���Q��p��5b�H�b�<�>]%z��ڊ߇J�ٞ���ř�W��o��!�`����,*��犺��_S��?a�J]��@����r�{\a9dd�:�J+`Q� ���+�Nh{q�/�SO*�X|G7��6����>%┘%�h2X��~�M����u�-�R������H���R��=""&?[��?�gJ��9+rR�����8	Εc�>�Zb�X��V=��`l�z����Wk\�'���ȣ��!��`��8oC�EI^A�q��,6�G�7P(.�^4TG����iV��WE�V.��3@�n�b.jo�)����7�X<,�҄=�����X[� �.�����[�#lI���HCtUP�������ID5d� �0G2,?�EM�W�h��O�Z��lBJ�'�3�s<KN5A�c`���|5��v��p��rJ����=�9�`���MI�^��Z���f��J��F��'bO~��v��X}}lN-�&y�h��^[Y~~���~E\���t59�]?В�.�Lk��{��TC
_�q�L7��"���M��qN7-;}��F\��~e*�Ƒ ���|A0�_��c�pJ��l<p�A���Ѷ�$ �`�yZ�Q<=���>�xw>��?�Ɯw�'~������D�Sp��N��	�6hh��;Y�z�-T�y�?�vsm�v#�pu�?�Í���G��~�γ��p�X[��c�^����4�i�:!�����S�����~�-f@�C9�3`����]� �D�%R榧f[���V��j���L8V|iwxR,rbq��̷�����B 0nP����I�?��9U�y�a01z�Ӓ��z��[l�uV��#b������x�Z�^�ց'��g�:ӧ౷*�I�ҜwtI��bB�kf=�ԳIIC�A[�/ �}��`���OH��U�r|� ��w�i�٩	8j�1���%���rL��-sl��e���b7�Q�0Ǘ��DsY�\��p�T�A���_!A�������b��5�Q�����w���Q����\_0���aB��[5���q�T���i,�ϙ�U��8 ��#x��d<�����5�46m�V���i��8�����F
<w�Co���k�K3��p��������+��Q����%�.�C!��x��0e�<)k4t���NkkBߵ{E"�ĭ� P^C�w�E9z��"��f�K�3g��bfl��;��|���;yB�~"Y������W� �צF�t�]\	�n�xY�K�5ғ"�,a�VV��zw�ʟ٦�".���K��`��_BC��{��&�𬇄���ڊ	�K����S��}|��Tɬ�[O:����ƍ���%�uYTې�A����
wU'u����L� Љ�RG{w^� fkao�?�~}��&���|����=���Z�_yY33����eմ����S��r� ���ԘM�Ų�tS�����K�6oٶTbU-i=F�3��� S@��8n:ϖ_��kh����b(��'���F�U��*���e�ä�{#�/SH�JXi���k�c������t�n���|����ɝ���m�]�|n$G���y���/����K|������$� ߏ <�)=����a.��]����]��)���o?Z̻v;�o�e�4s��@��u�< �͙X�Fo����qm��|�<'�x�]�l�J�'���N�hڄ����3w�w�u�{yÅ���Gx�ra�e��pdn�5��W��.P��5$E�ik��p�SҤ�S��h�7�����|�;m���:H�cA�}>u�7/�0�_��j�ck=�`�l<��&U��(�M+�y]O��ش���PxK�.&|Ϛc����
���[f��'�c�c7?ui��:�&1��b�(�������$��E���ծ��rY�{��^��,�*��`�Y�ѹwk<�8̷&���_]*���ռ���s�٦�����e�櫃�g���{�o�v>R�����`C=�PRi.#3����c�9M�Eɩ|>��ᝇ? G�@��T�WEi͈f�>������a�ư�9�C�;V���'4��L����˅ؿ;���*X��j4S}�O������d��۰�l�����R� f� ��S��Jj�n��÷3�Lml�`&�4������ߍo�lB��X�d��m=`�Q�IcQ�w�U����&��Ϯ�o�+ ���@!�_{�m�ׁ�s9�d�K��+}�@�9й���(J+IA*VH�>Uj�Ι�[��8�dyݸ��q|YO{���S���_T<Ħ���q��n�	L��ca�Rڽ\3!Wj0ٱ|Ay;�������~+C��/�;�"kDsoe�I��i^^�*i`P�s��/$䭄	�����CC�g|fz�#���\�^6WKm�Ɯ���!�����vo�b通c�m
إ��1����9��z��~�>/����HH������L�|Sץ~Vw-�ھ�;A-˓�πm�y�==is뒞ts�>�\Fg�ycgi�8"o� Im��%f��c���}�,.��~uɐ�wR���da�_5БۡE�e.�p<݅El��8����@X��@Ś}��(�����݀���� �h��R���.���M<%�	 �"l��l��_�:%���[����/� ��f.�3��\�����t�􉓃�VϜ"��og�םn�Gd��d<�n_hZ��3q�o���5V�{!�͜/:華��c�ˊ�x2i��_��/~�)�J�RD|�Y y�!H�-�xQ3"���Sް��e�%�C��#�@ca��H�UaR�t&�|�=��a0�W���������Ba���)�W��\�EJ��=��M�G��׭5�����	g~�T��:��N�bm�؝���hnHP~�5We��К+j+��`=:!�i�q&Ś�Nr����ɀ�".b֕iT(}���aًI�ؐG��E�T���<�4�9�P9�9AC�k�v����?�]\S���`�4�I���%9�qVa�{:S+�u���%+}��֑�9�s�|]��,�M�RiE^�/O]���Y�l-݋:m�q|gÕi���y����L������5������9����a��^�;�C^��I	F�����]�@�"�y*Vl=�gc��T��U
|���y���ѧ���'�/�(��8Iq��2-�B��8����1�bDS�n�F�j���Ǐ{�p�^��Y�+���kݩ��t��&<�|Pn��ShI;[��\��\c���>�fX�~քo?�?��M��dQ��|�A�-J���Qj�B�d�-�H<? F1��c�?�U%{u�9x�'B���XSe��偟�}���=�#3n �MFV�R���|�?5~p�y�5�C�	"�{Dٚ���TR��vq:sa��l���D�=n��D��N����B��K���?��-�.�4��Y��le�]��~���Ϭ+�3F����y� �0g5�;���:���o?޹����:-xJojC�L�<���ǫW���.T� �BpC��o�c��~ׁcr��$+J��c|�묙/�3P����Q���b&�I���-ɒ�bS�%�B&lzWhh�#��~D6�$_�Y�s�����[`Gꋵ I⋍a�W��UUZ�NL�-x����.����49��˯�#�;4xc�U�!��0}�T��C냃�x��psL���7FJ`�����c�����b$�Rbg���5;fN��i��և_��ܹ�}�=�K#0����������QHE���1HB Pq`�M�����K!R=��*+qME��N�Ȉ`B2@ؖ*k��
�`X�!��r���at�mTh�� 
��;��8��o��q�F�S��6�k�#˾�i�?��ȑ��!i�ɀ� ��|����bW���q/I��s>�x�f����-j-�{�������RK/hh�e<$K���-]�\k�ކ����{�u��@W:����SO��čl�:�v�֚��5������70,N'acW4��^p=6�=w��\O��"s]bUѲ�46~���N ���N�����Z��������k�f�%���v����d@�i�#^g�'�G���{	?��<�Cokt�|�\�`�NJ��w�{�����>�Y!,��c#�'i2(QGI�FG�#��7W$�W}v)�-;`��d<�8��__E[!�N�&���Z mL�Y�ε;� d0����)�7�?�u �����ą|�`��}��"�Kc�o;	5w��~���	�,;��^��d��ia���?q���i8^�Jw�<o��bV��@�&�`�0є{r�5GʿZZ��):A+j��%��>A�Ny9��_/u�I�10��8�
*G�e�We�5��uR*@�����&ðt���9 �c����(�S�`O�.6���-�wP*M�Ħ��ƌ_����&��e��C�������e��x������C̘(��U�	���N���9��揑����D��w�n,N<Mu��A�O��B�Qw��>&��#_'G�|z-5��ԕ_���@�ƻ�-"	��$<����)�Zj�VqT�>�N��ğ��F'�"	���.��m����#�o׫��
���J���7"�%P��X�u��x�eH��܊����0��:7��.�o��Yv���e�C=��g�X{�,���@��B��Ǧ|�� U8�i��1baܫԨ�4�<4���+L���R.t������8�b��%�����&�a7���7b�� ͇~����?�����Pw���h��i�����K+�X�^Գ��˰���d���z�l��Ma�t������<�g�hC��"�:�A/�S���D���	:�O1�+Ko;Z%�@r�������d2�o��|/,���,���݂��� �ww��]���lr���ުo
�؂}�g���93=�y�����Ѯ�OO{�5e��d�O�{?U��#d!M��^���;�
��x��@"	�|G~�h�m���ɢ�tV����Y�� �(Ek�n8�o�8\�N[�7������@1�>�
ΛG���A�oX�D^�n�bz��Y���T� ��n�"(���8ť���1�%-�2�k��V@�ݚ��3����!&3�j+[]��>��`[�BB�4}�[�1�ph��v� P�E{t���Pq~]Ȭ�ay4���ₔZ5K��`�KJ(��E;�g[�D[��Ɍ]�����|�Zߒ��XV�:���9���T�>��|�G�z޽��A��zz~�yy�}���%�|�>�W���!}*; �tPnpa�iO	_��+[E�3^b\���O`�28�~��Q�U ���-�������Zi����^N~P�g=��81���L���6/��AK�5Dv�з.�t��!�'�kZ�����k�`�}ԔЁ�`�����&`�^L�&��]�~SUu��P`�l����~�.M�P���]�\��;r��7�����M��E�Kv��	�}���wnC,���L����UW�u�����*3m��le ��k�U�Ip�>���N��ʑ��8��.�;3�C��2<�{z��JO[ �4�'�9u�<�1�tVY/??V��
�pN�Q��||Xw/`�~uR'�<$��:	S���Y�Bk&np$e{'��07{ACCo�QXVX�UW s�>�F��ǚ๒W�֑�����1 Kj�	�.�g\m���&�|[=5��Qƚ������W�~�6�su2�V�����Q-���ä!#�p{8�|[1z���P	B���G:b˶��U~a�^3s>���G�U؉6�[&��,_�\�� �T�k�)�Ud���y�ߒ6s�[T,1q�=)<������r8:V}�ʅ�X�}e���Z�P{�ۼ�9=S����M����)�90'��E�=�֬��T�f]�|�b�B��bX¥ivϵ�ys>�v!��Z,4V�� �%����!��U2�p�9���C�y,I�ȫ�2�ꭹ�ba uh�(�P(= !�[@Ķ-c�@��1�}h�q�ѐ�qؖ㣕<&�nbO5w�C6�B�ׇ'!Kي������|*���m'���D �i�E�*��I�U��K7�����BF��]�	��+1����o!D�I	T����ꈤY��R�Am)�`(�K�w�<a���� �~��(�T"�"��+���/\ D$�ctu��G����.o����?��Gș�]+O�A�-�����wݒ��[�0�{�&��6��d��ny�C��r�|k��u��gk�
�k�nܻ�N��|�������Gx���E�J�*C��c����N����I�D>�W u9S���u9<\yw�$����bzY.N �}R���D���<��u�/z��	�{�vFeH�EJ�B"�,�*���<�ҧt�4n������a����'��TO�J�7��c�
�j�����>��B��a]�fbye���c5x�5z���w�_U�g��@|���9���� ������Ѥ�,�1�� 
L%��Z.�?�D�E;$p/��D���к5��x��C�tw>۷� �Tg$$N���<>4�8*��up
�f(g�B��j���XG-
���+Iƛ'k�Q#ëk�����z�,�+Le٭� cS�1i0��v�a�t�+�W~��dՑ/+�?W�;�*_l���Psm9�����;@2�����6(0�]	Da���L�!���[ ��4��
�N����[j��RI�_�y<�k�c��/m<���5ȭ���YG]ѥB_�C��|���B������e�(n��=��\"���V��z$x��	�tx�5�G�q7�H���7�����J�x�(n��lx� =�s>����MFg��Oâƻ�����J��u�V�N��d������J��Z�+�3�W��U�>�C�F���Ga�Q�r�)��&�1���s��6�/��$_Ȉ���쇎����U��˦|c�b{���?��[��}`sK�G����_���-��6:��>�R<���<<�&�/��N��d�b��N6_�@X8�F4{9O�,]�Wk|G����	��v@�f�<�li�Ū �$x?*����֑�� �ZԻDNga3#��H*� ���f������Q�#��<��yHW��7q��+����l� �?�'���MJ ��ې��Zp�J����o��?��P���qy�h���S��5ٚZ'��ҭ�E���P�p�[F��g����ҝ��E�D<�UM������Y��y��6T�0��e�To�y���/����8x�̅�ݟ˅Y��՗�G�����k�4\��b�\ W��v[DBgN}�I�#^��_bpM<v��w��x��~��+�7ф��%+�����~AU�9�M��vsі 7�)D�̯C��u����d�Z�H�S��8��d����ڽ�q��\���d"Ս�u��Ͳ�=�1����� ��Z��vt������'c�	&y}|��5���h�U��T�7����}kB����w�n�Z�{��#�����Z.['9:ݻ�.N�;	�p��~���Ud���#|�py;�~��������j�8���"w�&`�s�2.��م��f4�]�	��n\ lmc�D
�R��wX>�+L2Cqi��}~Y����f^���f*��X��:�r}�z����U�/�ȳ�^G��H7n<oF�����Կ}.Ol��Řu�7W�z��7����O�RA�\r9ArHI�cZ��R�'T�Tm�I~P�_v��6��.d&��/�0~����2��)eԔ���H\����������O_"�8�|$��L�a�z���	����DY׋�e@ξv䭷�9�Ϣ��*��i����~�{�4;���R���1�������[L��(��Z��O�������t!�oض�t>�\��'��m���+�.��r̆M�̱]�����ep�[�������n4һ��=�!���=��� H~u�h�ӗ�+Gۈ��C�[���q�ep_��'k���7��(�C��r[k�_�^@B����,}r��f�H��L�/gE�R�$}��Pr�~&��j������Ǟ�8����7�������[yL��(Bo�XT������9�c����v�.�|!��n=��Z������x���T˛O����&��Ķ��� Fh�;mgi��9�b�te�N���$9�է�k�k�2s��w�D�6`|�g�2_�k�;��ƛ�d��hw�5*lB~p�p�XҲtF� ��کQtѪ�x�p�X�v
}>jM�҃U��4p|!l�XE�Eδ!�=TM(��F���#��}5�:|A��X��MhB-��7��_�]����#Q�d�c��|6��"q�,�MP��L��b?��(}�n�`��m䳞U�����%�Z�15ɦ�$W���2Z���=碾`%�㣛�;utk�}���].��/�5Z���]���J�*�/�֎n�bX�5�an�_Zc2K���\�xm꺯�+G=K�h��g=Q�	�?�`
�4��Y�*���	��u�>�<�
���x��t�fj��N̊eiz�ޜ(ע��k��s�.40��n'�L@y�k��)/H����^r���.�"������A"5���r��%Y��Z���G�t�s���;F��sV�X�vX  ����(}1N)�6Vv��O�*
p�x��2���MM��H�tb� \=+-�)dM9��b(��}TK7��w�t�i';�[+��X|�w�m�|pO����7��E=��z>��l�sYr�
�q?� �Z��[Z�mY���-�� �+�N8������KT�VY�dJY�z�&���A��3���z]������ث�׶���G�oDewVv�YTYZf��:o��^y�Mil�����g (-p��z���Y���9��;�a�wPőtW�)RN����j�M��E��ͪl�����~2k٫eQ������`��ee�#kg����Q���fX!68aj��&ܐDK�ޱ�xn�_y�ߧc�w3���V���4Q����Y��Y��=��y��:7q���������J�
��D� � 5��7l���C��cym��\�r�#��d�e>�f�yG��Ωe��_M��[-%��+�ْ�䞇�~�XF���4Co����SM��i����ˌ釦���Ԏw�b�Q�禬X/�rw��;ND�a��M?���K�EY#ʤ�D���>!|�$��ŭ�WS3ٰ{$�=-:��S��(<H˪��zJ"�jٜqޙ��͕�h�X�c��ԙ�G��p���V��� �F�g#69��������[�הi"�{e�i�#��[�Ӎ�e�x�U��O��s\:Ie�B���̕&�'(h�EǗ��u�C[=��.��3���Ɍ���i(̅i�H���s{n�����E�S4�$�o�Vc	�
� �y�R��#J����x�41z�G��w�Xmu�߁�;k�{e��&�Nd.����g�E/H��H�}sK���S~t��*��y��am����=��y��ߙ���4�nR��h�ImdP���Q�dߕ��}�����͛θ2����˘���xM�bϨ�����=�Ǿ���2�&Q� B9|.#2��-것�4�4�� �P���ԇ$U�=^d)�a�o����	=1 ��;�'���d��>��Vy�v5�~�����%���9��!|��Z.�W}��j�.7�%�?������0
̫n^�I���R1��K�so��m�$�y�4aÓ�`�x=�Nec�p��9t���0~fv*|�:���n�)S�ujQ��h�j��o�ۼHq~��2��S���X�j�cJ�.�x���dLso����݂��b
�ڡ��l�S6C�Yt���KM}C�ք�t4�|��|�H��m������]?1S��Nj��K�Ô 2�B���ڳ���A⁮*��<%;*�T�fsU�
G-]�)�[�|���i�2�h�H!YZ$�b�O`����+��5II��~s�xhX�؈/m(�BiVU��L(�ڳ��̒�pt������g[@��6'N�f��)����]�,�3�K8�NP�ڵJp�#�o?��������⋋�%m��37��4���.D�{�f^z��X1��,�"��ӧ�̝dǀ#���Ha����cKZ~�l�Pu�o�mN�!��<�E��HP�_��jw��|� ��}���v듛��1�5@��M����%t;�'/�2v�%�r���n� x�$C��D� O?;�Z�n<���
����s��C�kנ9N��>e���oy%&�����i�D�1��?00
�������i�D��b��^����Vj[�)V�L���mzѭg�Bk+#e ��\]��'�39����|Ɖ�P��L!�	�nh��:�ѝ�aA���(�<t�������V���	����",�Dh�u�M�IP ��|ʛ��>q3bw�o��$g;���_J��&v7�C1�G�-��F�|�:�3["�Oޤ��nPc�]���\�|���?���k#���<���p*�V��xY���k����~6��D3����C\����f��y�ܣ�B-�&�H�m0�|NI��k�a-�׻N�� ���_�Z�b\��|=��`>MǷ��1T�:C�K�>����f.�;/<D�\ҟK�D,]�R�?��}�`9<{�I�D�4;��?zG
�}e@�<�|�Y�̛��){�$�F�8���]un2��ӯ�(�y� C��ö��V�xnr��y���g��7mv���^Q�kh&>�ũ��7�%�b����g��$�{�u�H���.�o����<�v ��,��ۏ��*?��Q|��z0h�6(�@����ǃ]�R�veA+�I�j�?I���϶��'����R�Ó����4��{D�@�]o�!r���˃9��(EhiE�A����{O��č�ީ��3Cd�n�Tl�*����D�Hof����7^>p+^_^��� �]��MV�}A�: 0�^��Ǚ�4+�YAM��=]c�+��S����Yf��:�.1cm�Y�j_p�_ߏ_^t����� �"�j����t����`���:F���~�'���#6)�]�ǧ�W5N�o�(s���/�鯥��%�����?߽e�t�FD���;FKK[�4]��e�"�C���^ӲO����"*䴯�N�ժl������I�����Ƹz���+L���҄�cTt�3�A��pߗ�>Ȟ^��j�������ձ*:�ƵnޓRc^���2��ò�����`F�F��E��y�a�Ȥv�]�G!\��w�<𤋪��_��V���!�f�ˑ���^wD��'��Ԩ�w�}=��ʙ�'�Hz�ϛ�U�w�|�Sũ��H�"%}��3/�(�|�}���kH=�"ά�mgw]�}�ܟd�^1o�c5��u�y� �Ⱦ^/474��� w��ĉ�ȥ>wiZ��T��ǥ�/�-2f݁_��
�x>rOO�W�8�O)�����;c��I���k���qK\x��غ'?�rCt;�;�lK�9����+�d��0Yk�Y/�G��&"�+7
���}s�冖�_��J��~�t�4�-��)���������v�{���L��~y��>���
�f�_�t���=� ؿ/17�LK	�D�f?����U�v7]I�Ȯ?�&.��O0������E1��,����>�I&ї�1�y�'��\�,�/��k��T#�lk�I7T��Β����@���=�X�/բ	���Q6�?�a�ݕ,�|G�9�Β���KB��,�|7GU/�LM�;�W��\�x��Ah��	��m+ná]��؍ī�8�K����.@e������U�a��D�{��?��M������PIpM�M������rO`	Q�7*�����ާ �����;����'G]��ӕ�����`��i��g4ŧ��\$�E�/����8{�ҫa�9 ��������� }�,M��:��!'����@�5_F�R%_�a�9�d^}���dy9�.ȎL?��*8�@��	��,�;jZ)K4���>a��x-$ߘ���ժ��#|[��Ah̕p���u�k5���,��(}�$���g٫�K/0�6��  ���́�� �ܮ)��~�=w��ߝ���iy"����~^^�X����������Ɗ>ΐV��̩���[3AQ�~�Q���2�m��;
Y�bc�2c?9��$�p<8k��4�,Df ��ݵ�H�Hޝ�j�_�� ܚf��QE�_#yO���P�_��G��BR�oS��o�Q h�fj�s�.��i�Jl�Cǹ󽣢�L�@F盫�vl�sC,���]����x��v�j��D�x�p7!�e0��@����IB+g%6��`�x��bR�2�����ՠ��*T�)��m^�P�ҾA��st�CTt���s
�~k�G�O�f�d��BU���{�>ʮ�M�ڪڇŖڨ��������Q�(�����rf>~~��ܕ9��Ⱥ9ܖtk��]329i���
�I�Z���\���S,����F����H��̷��l8�+w]��d\Ha��9^KZx�'U���ݜ��(��N���i@��>��E=؎ꅗo�� ��뵺�����г�~6k���檸�}լ�'�%F^#r�������:�@��e����T��N@��O�e�u���m���=ݎ�6�oJ�wؗ�r4ȩs|����4�@[F�BG�IZdM���-�>���q�	�D�o�ASt��s�q���V�SE[?0�*~��L��m�ܢܩ(Ԕnrb��i��yn3�a����V�y�f94Z!ڟ8\�_)R���K�?�rV�{$�N�;������v���}G�h�`��h\����'�uFB�r��ٴ� �b����}�9����ܰs�p��š��]�ӷZH>-&�叓�����^�R���6<�A��'�9o���S�=�A��i?|��>I�]��M���sTC�b������h�y�@���?���
��0��ic�_�k��u��'x5�w ��iʅ�J�	9R��!,�������o��w(����(���w}����7���������EM9^��FFu�n��،������VΖ#�E~2��Xj�d�I��������>�FnjpS�Y�MMt1�:�V&�붟�%��~��B�0����m�*e��t؆���/��ǒm����O�x��a�6�|&-�����P����BK�9]����*��O`�%a/$�z�����w�;��՘�ʗ6���T԰�R�~��ęH%�Ɓ���}v�o�މ�|����ʵ�'cs<�/ia���w��DE�V�%\�1����GY!�)�Xy�'�1s�xݣ��)��c�a�)TG�?��������^Óv5�,ڊވ��M���~:���/7F��D��w֋�B�~�2ќ�0�%��3�zG����v\����M�Ӊ7��'�D���:��Zs-r�ŀ+�WV��S�(�79�<�pd���[��oRT!��+I���~ L��T��,Z�%�dv!�zF�{G���ͼ;w3�f���q�Ta��4�U�������e���"���c��^�Õi#���]ua%�iW��'O�yg$<����w��_�6w�����h�V�,�g��M���2�y/{���h���c^?�~��qM��:<�����3Z�u]�*7`��~� ��bX�T���8u��UZ�g��D�q�d�#��jG��dѴ�˾����H����o�#�[�4�k�e�x4F[�@B2`������z�_��ߦ�ԟ�]{��לrdZ_��T��6���qN����{�A���=�aÉ����Ʈ#]��:�,���܏S�jw��u�7/�y���]H�Z�S��2�G�a)>��A�.Y��*!�����}��c,�+~QX����-��"�@<��;��g�0(�jD����=���Lr�J|�7���}�k����w��L�r3A�RTJ�gps��:� Ԣ�(M�����|ѐ���j ��x�/�����h�?Ѐ|�������H���~��L[�TS5;��T�D-%�I���2�OU^�N�۽rKT�-��,ݥ=�����C4����:B�ߒ�m�P�Β<��M�[|�"��X.�9;�l	y�
��+���Oh(���s
>�˿X��_�J6x9@f�!AVMU^Z�C���ꄕn+L<���a�����+��e��݄(z�����f�, �����8��a���wR��k�8|89[T�h$"���Da�Y������;w{e�h����E#M��Ӎ4~����<S��$^���G��:f̧ݲ۱�1]���{E.7�I��c������cN��[aw��a������e���Y��i�z$�v���fok�r�ˑ\�َ8�I��5��y���nY#���������ʷ��ED�5�����[�3-(�?�I(��I��W.$���f �S�ƾ��:��q$�j<��#�����v�ˤ/P�؁�R���q�����8��o�X��!js¥z�����͜8��ɭ0���"����O�Wdx��Eɲ I�˱p���:�T������9�?��i�T�[-D���>�p�����y�9�K"k�������Su�)�ۏ��	�JJbKS�b/%8��0qS֍Mt�y�k��Tfڸ�"��*i_EJ��#%$��ߦ��J�����$�x�ᘽ�5[;��x�%,�)���0������Nֆ+��j݄��Q)��:S��gٽ'*�*�2S(��W��ǐ@���`�'`���<�QIo�
�@��4�P�w�.L�o.7��b�X��9�0;�u���Kz�UZ�'�y*�D>�����������<�2*x���|���S��ߗw���-x|�(�8�������5uF~�i���ф��Hw�O�z��9ݣ�YXۺa!X22M�كJ�z�fǊ��	�(ǻA=r>��1d^�(뇓��^���,i�Em�	W S
9*v/P[��ex}C�C�>м��@D�x�Dm��GS���u�7_����1�I��v�i^&!����هU�R�����>��zu������d��=E �S�s2?�Q����]3��G;��R����҃�II̧b��g%v�v���Z�{��������j��K�T�l����c���� 4{y$��%�X
aa���C6��2V�k� �Wy�z�}E�I���(���cb�IႨ8�u�|����Q��w�{��e�n��mSG���˕��OҒѣoK���gf��3KR��&��g\����r�Z�W8[�F�D�Z;�G���~t�C�-�qTZyxtB�q/<��Zf�l���0��E@�o��VB���ݶ.r�L����(�۠����]a�9�~Wir�k�Eޱ��;�Wr*���7��v0�P^v���H���~^�G:�潍�5�F�uՕJz���'�������Q���)s�XL����F�reͯ`��J:�sڕ��_�T�5
D�O;��±�o�_��quY%���0,H����h�f�D<$�a���\��8���n��TB�r�ۦ��C��_
a� HX=�3���]�̟�͖��C��7�_Z�:Hd���f3o�~Р����_�)Q�Ka�O�d�d1�b�_9�$��^����{u��b~D�<j��վ�	r�-����W\h�4}�]��qY�0qe1ќ4�����zD����fe���U-�A����v����8��6����&
���!��ȷ�k���v�G/w�4%�Q鲫-��ݝ���E.n�AcTt9|��=Fp؛�h21!ٖk���� ;X4�׮���ݮ��N�F��z.6�eԳ-�&�@j��ׁy�n�鯺b�"yR�ڠ�g�C��3N�؂̖��:��F�G�CDK�ԡ�l�����66v����E�@p�Z:NԐ��`Ֆu�ʃ��r�ضL�d6����oq��f�'�'�L����4��Z��5�B,��j������	�Z�c�ɫ�#A1�a6�?9Q޻l�1c	H����FY`��#�����W��4;|� YP�D��If|O�9�"��`�=�d�^d$ �0�M5Vf��0�D��f+G=]��Ʌ�hK����m[����frѶ� ��6Od� f���P]��+Χ�a��fS��SU��֌
nZ�UAMի�H�(��?�4�/����z�.7]:�ndO)��37���x�J�j��%�QGd���b�wć�۽η�׆o��<V���m4+�ȡ��5-.��q���]���S P�Eߟ/�������* ��U����5`kh����n4~գ�f�7lf|�{)&�r�������_#��S��M�V�y����ӾZZ� C��d�Iù�T_W$�oō�c�h���=���/�&*���H����mS�SƜ�ZBS���cVˇ,5��E�*[[��w����_��}V��#����[�n
}�[4(����K���e��w���C��@�8V�l[5��H᠚�Dh�wǣ��M!��0qsG��A��JX�{��������m��z��6u`��'Dq��ޖT�T�����8e�����nI�9�svWni,�����ܹOT�֝��ݏ�<5�	��s����lt�ؒ(�6ya�ۈV��M7ݩW@n{+! �M��(#��y�?�jO���hc~�� gaAk�̯����Yˎ/@1A���,�@ ��Q\�Xu���Y#�i{�bau���^tg��te�˄�E��G���?���Q�,�[8�.����f��?��E�5�xa��N��<�H�y�P�N\����7�����c�Rl{���#�v�9�|���@0fV��(2�����(]!�����DՈ��u�.mj�p���v?��e����T
z c��M6�<�.+�3� 0��m�1�����:C=	��~�X$'_3+�=,O��Z��|���c,�����mz��m�4b�T4>{Y������+=bN��c
�ARc����)5äƦ�eL�Z��?V:�������ܮm6��8����Z�ݪ��3��z�����`����k�2�A�,&�L^7����M��_��B�?7ZqsĒ;S֧E\�e�$l�Ǌq3\��1�JM��l|��b&���&� �w�� ��R�I�e��)Q�s0��ʁ�ʌ�����x�Z!��n���߆��d��.���}~e$����-b_�� ��,���%�[^�]������H70VV����]4Z�A���OZLVR�ud��$�P��u�V�?�11��� 7�`6��!xY!ts�/6sxX�g�d����,/R�=��EqZ��泮�[L�'��
*���ͤi��M���T�	4k+��\ֆ��SԄ<�[ll���1�@�N��љ��wgW�M5�� �z:m𞤱ϖʒ5*�z	>&x�=0��I�,�ܵj+5|�2!b���uin6 $��I��Ad�q�dGҮT�%/��P�T�M;e��E���l�y+2�=	n����������%6�(�W ڿ+�����s=���#J��'aȝWfJ�)c`�gCt���V��Ǡ30Q-�S���Cs�~H�?��|fL��	�� {���<~�9�}݃~Ck*is��o�L��{��^���,m����x��!�8[~������]JZԸ!����8�����6Z��|ԥi��O�mCfWwa����6��� =n�\�կQ�5��P����LX�1+9�4q���O�xc�Q7�C�PS�E��صe4x��Y�q��
4Ƀ�FjY�>�C<�a)�5��l폢%*ʵ;�������W�3l\$dX �(��B�x/��������><��0��j��_�n��J���$M�fv����?�J(�:~��w\:b�~'2�#SLE�8x@�	^4�������)9O�v�?��ЯT=B�pwK�YA���VA1�o���8]�!U���\�@�:o��p�{^���q�eҕcR	P?��jM���N���F�����X����SBgޝ�;��a'���}�Z]	
 �c��H�;8��T$�ڕ�}�%��_�^��>��T�K��dE-���~�O	�6�	���V<?w��ҕ--a�� #�Dd2��9��}(9 k�n�MRj�.�iL���ޝ�D��S�t{qmؠo�Ƥ7⃃�+{JE�`@غ�פI�T�����
��w����Q@�m��'�a�X���\]BM�w�:�]Y_y�A�R�r��t��a�@7�=���p�e�*��_4?��A��t �b-�F�J�i�5��}S��"���6�����w�qN:9mL�Xy�&ZO}��h�L9P\(,��Ǎ�1mL�?�j�"mǑ
]zg�þ��P��|�\�p�����S��%*��I�N��'��;>��K>'c�K�el���x:�D�D�^\Wt%R"�O����`�b!����$
��� N{��G��J@��h"/<>%��ſB�w�C��\�%*v�?�����{�X�6e%M;D����ܺ��;q�3-�Kf�(?�{����͞��⠒(�Q���Ϩ��&��۫"Jy���׃R���^���M�Q;�'���v���� z����Ҕ�d�D��
�P�/M��<OJ���a�[�U����B����b�?�w1�23mTp�z��T����Y�0լM�,k� ��h�z�nD	v�K怐|k�$�揨�.iw�0�3������w��`�AP�A�%M��8RT��E]���U�RD��ܰI�no,�g�����moܖ�f������~$��Rs"�V�m�0�S��B&	c�#^�@]��G�Y�3K�}���v��
g�-�C�Mt�[2>lB��\a���P��jC !5��::����g%1�'/cW?T[9}�$噋r�p�X�o�,�ۺ�4�O���G27[c�Y��Sk^Mͫ��($?�H$H�G��СA��/ҳ�p�/2a�0����e�y,�\,��<���QH��NR3�JM�Yx����1�?!#E+��h�;	�;9�e	�U�����tW��w�&[n��bQ��$|0^Q.�f�әG۩]1׭��ؘZ��T܄��!��v�1���$���+�	�w�����I:����� �+�1��{b��Oon�ß?�ͮ�M�����>l��;����5�Y�Jl��t��u5������6�X�֣o�[y�gQ����'�!}k���f�XZ>\��s̠Ҟ���H����+B"��4B��B�C���mDF?���K�O�ܟ��[��\�����	�V�HS����]��i�́�T��!��$b��cR�����)C:GLܗ��b���!⸵����%���t���R�XҦ>�8a� Z���� ����\K���/�K�)'���T��Z�1Ŋ��?�
�K������ؙ��%@$ɗ�)����8���1�F.�@�dJ��B��q��~yY(�q�Ĥ��h�ɴH��h�;}��6V� E �����GP�����}��˂!���KO�u(v��sT��=}�3x�g��O�:�/u�B�������l=w	Jڸ�|��A	F����@��4��`]ZvI���R�+������4�������b�P%7%-U_�t�޹V���t!���Ak㒦z�&��.H��.���v���5��{y_u���B��>��*-ldR�GD��� ��-�P�E��4������2��/�(�A�y7vd��%X�����cfއ��]B)�?��?y�����,b6_��W�Z^�!�X�w���+� X����0!m���ܴHϭ����������r�Ҋ3# p#{T�'W��7"�:��l]�3�?�p�c�X�ԏ����W(�@����s�RC����g��K�<��-1SU�'����~�3\�����s-��ō*`�?� �>:!��綕u#Ţ�; �$R�YW�iY��.vt�	f�C�u^�&����A�$����(xߦ�?�$]�"+�	�o�
���^�2�J
{
@n
zRl�����.7�<}�����*�Z��N�(3c��𺪊;A2�����#$�>���F�IQ�DR��\����h��3�-W�ag/�eT\׊���=m#C�LpK��oYg(]��|\J��,�x���$'z�x��z{�P^m.0��w%=��tN3ڿ�fA��OKM]��P)k�u!j@���6!�m�ȷ�pu>Vj����7����bh�KnD��!�&Nw ��K,l�'Xgc�oz �,�{���|Bϗ��yY�%�{�%չ����I�Zs�K�y���?���)F�f��q`�`�d��,	��#�KBL0iԂ�mg������.ǈD�6�1iN�+/���Wy�5��9Hj��@ �M�?�<�z��f��� ^o��&I4��R%���̦�g:��CGQ)��>�2�b����1�k�ͫm%����U3!eG�/�l%� �A�9��GlB�6��G�������J�7ǥ	3�"��D)���O��iA�����i�j+��O F��I���:��IQAP��e.W��y��Q�U��+����Z@����Q����ijֱ�-�h�Ѱ
WX��ېƈ��u��K��v�cI4�2��*��^��ĭ*yG��
��_0:*�a*���V8��
�������g����t�ˁoue���M�V�S\�CJ���ظ1��s*ݤX?��_�?��Fa+�1�SȰ�"?d�b�y�pt�
PZ�XA��*i��'ɼ0회�Oݛ���~,|��1�[+P_:�M�1�L,���HK� r-���/VS����� ���d[�ufW���K��J@��5���C: ���-W��dL=�J��������\�a@-nS�D3[Ι��o��{<:�2��oqV_���!���"Tb0��B���!zN�Z���w�,�?Z��T�S% �vv5[G�|Z���gr�������ݝ�ly"Ф�*M�Ǣ���]{:�����|���#�L�H�	�kv���^� ��#�S��c��T(���P|A :B��u� �F��xUȲյ��Aܢ-fϫac���+?�ճ��P�vv�~+����,߿"�ѡ1Jm{4�i.[_l�fG��~��� �w�+��~ ��U{��xd��7������;a�z��$���>#�+��ġ>�I�`�\���^����y��܀r� fk�MB� �j[�Y!���4�"���>�7��1�������4�"[��mv�W�|��I�f
�5M��S�l�x ��ZwBj�`C4��\TX_Ml�'�e�U�_����Χ,��S�(ݙD�m����	�V��}�Z���w�� $��s.z�:���%1b;��<�$�PM��'ur��z������/�����h���R�]�
������i�ޏI��,�ח4��J�T�C����ϧhF��K�׎����B��2�z�o2�z3-�L�0NL���EďG�n�IuNr*�*���=�;Vf6/��M7�\n�K�~;+���F��L� �.)�7�� ����
Z8�%�H� 8�-8�c�����?��-P�OMd�W2sY�Fbk������'��.31� � �b\�x�
�T�*�ʡ�.�����S2�E`�!ﴄ�䞞� �2l�"&��@J_/GrJ0-ψJaک�\� X�_��0N�l�Q���$��E��'o��З���]/���7�X��)����š˯��ʁry�����w�"��U��R EGE���+��EB�w���?�2��`�ָ�Ip�@��'��o���4�ww��v�s�s�ny�g�jջ��G$ю�$�(ǅ�Rp�?���tZ7_�M\CP��m�;�	�`?ln�GEF�Vf����UXX��ˬǪ ��>|��s��뇖K��ܚ����G[���̾�	#=�,}nb��X���>��%Ʀ6�c���,�=���Q�Y�$�F��!瞆��8���z0QF&K�V`JGQ`��(�u|2z�x�
�#�w���#����'V�:���W3#ZXΣq�8��ˊ��v�L��#&��Q!�x��p~���)�/n�+��ݖ�/ng�d���`7��@����i"N�i7�����;��@��^�%3��Z!`,[������&���g}g9�	�Dl����X��2F�^r�j���g��#���' ��w*<����'�U��M�pz��Gg��+�ab���	"J w��cB@��3P��E�~�Qo��}�{��s$|��MZ��1B�+�:J�#(W,4�U�.	� *?E5�Я���B�FR����R[���>�k� �z�;g� ���7������e��/�K�Ќ�$z����$��/�T��r�k�mu9�=a�5�q���������#Di���Z덄_�P��Kwe�����i�Q�t���s}�O�_���&�
�yt��v��=��0\��Ԗe#EI{�0��W^c�{$E��7�_UN�s\e7yef��w�k���,�����7�-�I!sw}���&��.���^�|��>��� F���l��ZTe�F����X��I�����
���Kl�%��Ƀ��S}��,~�����6`�Z�N�� /�����䃕�M�N:�9NF��q?�~{�v�o�P��G�	���$b������ޠ����A��{/���DԮ��+P	л��ǯ���|'�N�U�Q��P����<��0��Ԙ+��	3Q��Yg�~���|�vb[�f�\H�P>����\�'��k&'>��*��\���A��Ή�`��[�w��q����g�d�E&O���b�����QN��F���H��gN�^ЇӅd��7�P�72kq�����w��@���/\�a��iVT��+2`���8���>�_�����}n��;U��խF�-�"�����}��,��K��۾k�e���c
%}��'�c)�}kL�Q:#�86J߻���;M�p�˾�G���a�&7���N}Ӯ��3���]������P27;���!q��?����y�:�V��chMTg6��~$"�W��n��8Iܾ�zylhaXkd��l�Ф~��론��E�+\l����_|� ����(]E�.D	�K٘=�E�I���A�	�?�߸X�mS�N,�w����QA���K�㭵��HL ����ZJ��"�Ր( KZ�nw����<2	��V	QzcS�݅�C�T�i��C'M�hܑV���a�㩚jo�2͖�R��m��-�{l+B҂�W@Z�H{S�W��i����zwdC���B�W������1髗*�O�?6&��-_0��ӈi��CJ�̟��	i�oH�Aۑ
Z_W���~"��+�P�V/�ɲ���]s󿒥ͧI��)��
�{k����c	o73~j�'!�(��۬�ޚM�l�nm+�J�/�L�JFM��Y5r|�om��7�ջ^+������j�kY��@�1۾�{����k��з�ؠ�k�NUd7Q�8=�o���2�|2� �k=��C��N%OR��]��&����!�mg�nL��KHsQ���K��K�Go�e=���e�ƹgU��xgs7�]���WS'b,�;"�����G���XB�q�C��R�s�ǲ�J/N�W+#O�qV"|��P���(�m�)~B	�|��4c�S/R�'Y�$ ؝S0;�֜+�MR����P'2{�x��)O"�]*�]DN�qi�Q+)�⣓õ��s��P\�'���
��&J����_�7�T�o��Y��?��R�$<(
2WjU��6�a�;+��"�I�M���ղ x���{��Nh*ǔ�\�F=�(ص:1���z|�B�D�7ű[��Z��x뒞����_3���D�΂���0������!�2�)/mV�`_�(���F"WS���A�o;��n�u���D�F���4�>ɓ���i����Y&fv�z�V��[���A�8p�e��P�e�m��Ɇ�M���J����Z)<!h��Vn{�6Q��m����ʢ���m}UΜek,վg���x��^��#�D�.+8��G��Fǰ��^�e�Ůk�tgv=i@9!C�)#�AXa(��E���J�t���14/�x����s�c�4�0�\�Ƿ���M�z�+� Ǽ]��f� ��w�r"c����%���S=��NOGh��ӄ��'����uʪ�?3o����d�d�~S�nb(����"�6�U��Y<ʪl�MW<Ҋ�"d��lV$��JN��"�h�/����X��]�����q  ��ɨ�QP1���Q���*<�>:f�X&����b���^���ϧ:q��?�,|4,��r$��.R9�[�U}ZR�-iT�����o���qw������<R��Г�e��k.fr��|��Hv���j�\o���Z�n��w��.����ړc���%./׽�(�׹���/�I��w�N{_���o���N�7��15�ױ�����'�0'sh�bz[֒k<Im���PCH��9�C:/�<]�F�G�[�k쌇�5�wf|��o���Uv6���U,�g��|�ɉ��E�"+p�b�3�CB����f�;:qB��8�8x����
 ����w��[�8L/hdv��|u��^Q����E�ΗϘ$�Ł����[{�L����ԙ~G��<QUwc1׃(����Ȑbs�IbbD��P�>�y9��G�m*�'#�J�I�yk�+/���d���n X���y�J��(G����a�Q�.X`24S!uzIN8lrNB~�%}��o�ӈ�B0"�� ��[�/ڏx��4He����gU�4�_j�Y�`��n�P+s��ѽ�_#�}
V7��&X���{
�N$O�>��cyCD�EQ+/}� �����)J�2������/�j����B�)���	���W)�
SG�o7������ي2��y���x@`�C�+��j���#f�)ը^�U�r�E�m��'��AN����u�.�|���1-�/]b�r/�[k�	j(�:`��=}&|9���oޙJdN��E����ۊ�5/��eG�io�ǽ��U ������O�������\�.��=��[����1��V��U�^������u�4dڵ(o�a����T�MTE�ʀ,����m�P#5�=˟x�h�N�AN'lM`�ý�r9v�_7b��fi,����^�e�z�n��[ 2˓v�Y��5�G�̋k��� ��RKˁ<��k˰��=n��]L!�ڙ��∻���+��1�D������D�J2Y�emʴpgH�R_u]�X~�%��c��[��K̊��N��앱k[0�)��)�[��!�X]E1HZ:݊ŷ�˴�T~
��e˧=������7���|P����rN��=}�y�2�b�{�
�'jŖ;~~A*����^�S,il���ˋj6�?}��_�%>�����e�Y�bz���؂� ]c
O݆�ȧ��X�c�4�Z��;aYC=�_�*���&^oT�J��%C�m����S�� /���Qy�}:�:���#��"�]�����&PUVzm�Tl�7vn�U�h<��e�apzP�km�$�o�cK�p���kS�-�uc[���;[1��D{m6�����g2S��\�K���E#�Rw���	<m���mT���'�ţ�B�m�Ϋ���}M�"���1��$��R�ܹ�^��c��\�/:���g�G���=e9��6_w�_v���&�{�Β��L���Ŏ)r�	b*0�z���@�s2�%?[Bd��P�XX]�bo#gc
��+��f���>�ϐc#���}'F�@������M<9�Z�.b �a>����8aٯDe7�����Lߍ��^DJ:����켮�g���݆��W���#�Cp�37��X����p�sRQ��!>n��8�zUm�7��^�Ȁ;4���Hŷ�{�0:ޖin'5�w��~��:%
+nw2����'�W)���H�u�Y$>7~ܹK9�q��p�{�&����!�x�U���f�oQ�",Ϫ�]��E�r���Ã��s� T��=���>�2O>ס�����iW�I��;��ދ2_;�_Θ�}m$�@���gT�Zs3�����ɛ�M^}��R��I�D�?����[n̼�����Nb�>�լU|�!�����Cx�b~���t�:� ��V2�B�-Y'�p2��T+�xb��ZVĿϺ��u</�K�r���.��ȹ#.{ bKQ\��uj���_���1�U,���g�����t��9;�I(zoB�r�X��7
�87��r:R�0K�Z����r��P����?j�VO�O��!%����(��?��(,XX�{[G!�Չ�,�D+yD����	b2c�c��e��O�R(�xuC���T��TJS���v�ҍ�x8�r��<S�e�����(|XL{?�}��5�U�ܶq�P�,}W��d���^Ճ���m>-�LwwX��p�tJ�Y�~�0�}�¹�Q�pc�9����ۧưx�*)iBS�Y2�~�Y�9%��zd���ǳ:C&��
9v���Fhu��<�ݨhM[[[��{��>�m5�螘��m:�}��3N�P'��ds��&�S�q�ÏnSw�E�V.�[*{��zN�>0����\�/��qHH�'0jo$�����?��^�lU͍&+b�Ai�|�d��x�-�M��q��-���_3�TR �y=��"Ȅa�
���4?A��E�8�+mCބ�?��=�줐� �ņӞ�H57����Tn��3��]��|���l��4����Fb�J�����/�@����`�6�3 ����mϟS��ك��	gÑ{�;aN�"E�f�#�	���d:S�e���u���[� ��c��R����]bz6^��F�"luE�[����?�iI�����>�8���><;���8���ח%gXRש�j�d?��|ص�YY�{��N�ٹ-|1�˩U���o�[/<ڄ��a��@���i6�ˍ�?�h�Z6U��S0�B��W���٣��K(��]]�n��c�Mɻ!E��&�OAĸ��.!��Zu܃'d�c�`��o<������w��W��͘�Ȩ��A�,����OBo�'CB����Gю%G˒���|��h���R,�mP]�K��F�DDx��[k3��
��OG���3�k����E�yՙ}��
��&��	I�E+�+Sw'�D�ۂ^jx��1ߓ5�H�1����gX%bNR+�0#�3�FN+�ұ7��B��{���Y���]z��Fs�4��� ň��ڸ{}�5_�S�����$F5��@�͑���s���J����p�ٯ.�&��<dՉ�E����1|�Q��cy��Y�0/�|�K�t �"��k���+�s�0tK��U�~;�������Y��w�^S�U<]I/�j6s��@�J�5����U�H��V2i�,Ui�7 6�;���k)�qƏ�w�B�g/.��ev�y���s�hm��4��D �_����ͭ�jdo��Z���z6��j&�BCV�<�����FE����46��R�t�S�U�$�������Q@7N%�(cZ���+�'��_�ԥ�1W��*�w������y��2�w�� ��H��2 ��6��v4�0�iU��3��5��lr�$��-���-8'5�w$=O�D&:�@��$�OD�=�zl���Qt̒hL���$}�=����Z�ή�PP���ਨ�� �k�4����'Fx	�bp�Q��K����#���3@WS�T��b��@��%��,]�8 i��1؏[L�-�|JG��ն�{��N3FTw�<��#�m+�,��p��-��J%Ǐx�g1^�Q�������&�r^���D�]o�.1�>s)��}Gm����D��C>m�ko��rw=����c���� ������qX�Y�i���U����l���<p������O}�0��ApF&��B���̹A�!h(����,��[g6���1]�������v;^���V"4�ߒ뿒l\�O0+����@��a�����s�Òe��Y��2(�t���{�#������D��4u� V�^�����/�e��7*G̈鱯q>ǖ�����~�|�����A�@j�!ꉋ�5O�S��D�-��W`J��PX�!�h�R�����C��O�b�'z��� Z�H���y ~�S����R�����y&I1���Ά}�2�8I*��XL�+r�#$��sXi-Uo=�A���˳V�v'c����_��=�A	�aA�M4��ӹb����"�*[�3����Y�t4_�/i�6���S?��"$"c�5]n14���{��b�?�"�G��0�+_�M�l>4	��о�%|z��c9�ܷsc(jǩ��.s��BۈA�#g$~o��FO�ZU��:4�6���j �w{�-{X���.Q�<g4����T�럁oe��^[�!E��6n�ּ��a�����K!���U��6����pq[�+k�\:.A2���9g�CA�F���K��HK�z�*	v��N�9��2Os.p�E����4~%��6�M���,I)�]��ry"�_�~��RQ��|jg���&�\�tB7��X��kx�IF��4U�����W~�;2Oz!%~�f��ar��kToc�$�tG3�#��2��K9�Ȓ��:���ŋ�YAZbb��/���ZN�����h��h�زp)�����[�PE���DpF�]���/���R���9��&?�d=�����u+�I|L���E5 - ��d�E������(π�p1�KL�*&.I��	EH�\.��Jy���F;L7/��q݅dB��2�榗�v`C�V����*���Rŉ~gZ���F˵��{��ݾ��]�p���#$z��)w/������f�zlp�F����}��x���QwmTr��y��W۫.��;��cj8o��������{�GwʅeXU���Ǌ�QτM?b��W�Dg��;STG�_��W(�����s�H4H	�\�y9�"�o*yI�P��ɢo�yQu;�61����6��璄�o��YƟw�������h�N�9�څxȴжL����q��7+6} �j��$���;�Ś����D�طk�̫m�ْ�mcK��z�9���Y-�Z)/����ɰ���exLt�7�������˷�t��G|A��w�˒�9	pH��l1K��3�������S���l�i�Y�ߔ��i�@xdwd)|�Z�j�<�����l��Ro#/��goT;�ɞ��d�P;9!\��.8�q�L`ֹm�_�����}�mli��L��ߝP2�y��=Z@�1���;&��J��wV��7����R��ڢ�r@QQ��7z���պ�����������$9~I��t�px������=Q�QW�A!A�%�x��o�5��;}��B?0"L�'����%�������Qu)�=vT�E�H��w���2!2�wݑ���A��3�Żvﰱ�@��Q��>W�W�ȭ3�}�����g�=<C7-t�6��t�r�ͪ5��z�/��fR%h��6����>Lj8pF�jg~�7 �m��E"��+^n���m��Ō�ɉ�
G.�K�=E��T_}2�P�Y�Q �a�6��aס+_�TE����������f]3y<����J����z����8y�qZ,cRr!��i�v�J�J�Θ�!�'��Z�!Gu�C�}�J#��I�M�L���\��N���)��ב��o�$	�CN�{���)�ׯ(�'Ÿ��3�/��<D�-��|�񑔣��U�G��B�ӊ�h�-��L��_�m�6����azr?���;�1�8:8fh��XA~O�^�B��3�r		"��g�-�7�]�����Py�Gw���K��4���(��S�����c`�ڵ.�١c9?��[OON;����Q������j�S�D��o�|8��W�F�=A<��o乮�d�/w��,31�i\��5�a7������:��L�z&o�B�b>��łpPqq�K%.ς+��Vd��w6n҆���X�Va8�����5�-��3Xor!�q�p:����eR�q�]�].;� (��$�����5���ɣG�鶢8��-���95X��"`h�r�醾6_�����J�I���E@��[cs������y���"L"Fv�z�.�FpZ�>�n7��b�|�4�S�@��. վ���4���l6tίΟ���ݑ��y�]陕�0�de�K���ȊA�'��+W�S�d4�O�t�og͕�t7ͳ\M�y�+^Y�h�	�k?Fb�p�Y��I�B�ߊΏ\P�Ԥt���+���\�%X,-E�kq��|���\��j��M��6&��d�6����B �:�o�����0Ȅ�(�� :�wAZ�OVkkgZ����9]V�_,���d:Ō�YT$�kCT��lq�f��q�/v'���D�>dar���D8��s�M��D��t~@2�A��ڿ�sC���|qx|Y�VIC�z:}G�!�f[��t[���y�l�h�(�v(N���1
�0�F����iDɭ�h3�7F#�������<����zҴ��h��(�99�9�Z���9qT�8j��`;$��kn�=&>���[�ױ��\�;"	U�~HQV墛"!���g�ao�϶I���,H~��e�e	��ӊ>DT:�
�J��P��Ӹ�������b�+�`��F\�N��2���u%���G5�-<�]��m��O���ʊ �l�C��n��cK����tJ��' �\c���VVq*e�ɼ��G�>��0�'��P�Z��~�O�������Ә��M��&�m�RsJ�$�]*]�j����;�
?��ؿ�$���2�m��]ߙ7ղ����2��֪*�.|�qY��cdf-���	�<g�'��j�,�n��ˢ���Y"0�B�~������C�]�CT�Q��C紌�N��i��G3��\��3��+|:/����>��r��L���Zm�?x���f:�p]�W�s="0�J�hw�����m-��k�t�o�s	���������>�C�
�YSOj#��mcy�:T L�m��\P���Q��Ct�~�Qi��X^�h$�Z��o�=a!{�E�r�rF�����,��&�T(��{	WD7��Sd��t*����>MxQ���G0�|y9(�	NE�Ca/���&j��蛞���w7X��V�V����q�Y4���+̑�GƟ����Be�t>w~&=O�9��y�����<���14�CFC��U�\40!Vs�R����k+�\��.�Q�۝H�7t����c{7 ��*;o@�n��	�7v�M˺Q������\CGR������Q��o�ͬ1d��.~&g����ڝ���:�����oH-��t�/ʜR
e��}����\�/�^)�۳��GBdd�?�-At�������Os�c�oL�&�Kڀ~I�4��n��\����$�z��Û\�!�~Qs�˺��Fރ�+��V�$�f�����* ��ylJpd�-��.��}�u:�RR[0�z/\{�5X�d�Q�|!��Ӕ�Dt��Ug��oA��0�@�i�cn{����M.y�Y��b`��[#��f�9E��Uf�C}� ��v4bR��=�5C���E܂U�k@��λԜ�jCFu�|`�pM��S�=λr����|��?{�>ψ��zutJ��ޗ�dg�ls�M�zħ;z6B��]���H����o���'�'�ٷ0����b�1�j����Z�N�ׂ�����Sg�NN<�1���w�ظ�I�zΟ׽I�oov@��2/R}��R~��T���1W~�pg#�d�p]Q<3����?�*D�G�iKϸ�H0��MԨF&�W�����ÿ�m�҅r�t'o��c��눾�)����?�+KÏ_7`0�@kn���dlK�����\���}�'�d��C��U�E��v���eƋ�!|�X�w�#�c��y+�9�Н$�B��(�S��� �s����j ܏�q��?`�
�է{���zR�-���:�(E�B�%��J�����?!A'''�	����뱃�*���'�E�.���O�9s�uҭ��vdHwR��Pac3�0����!��5��M�Ƹa�Z�����_�c�(b㼲����J��?T��?�ZA��n��o�=���%��
r��)&�}d\���(��̷�����g\�t|��K�%�c��!��j5��͞�L��T��[�Y^U��2����x8�J�Pնv^����d�*�$�-ޑ1׹v�E�Oy�����o�L��R�s�������!��
C+�t1�73_y��$��������\R�t��cK��o�9G�sc�B�T���E���pR�x����dt?X>]x�ͬQ�I'J��XQ�B�Oe��0�g�!�Kٴ��as���z@4Ӗ����X����[Y����f ����D\<�,@�,�w�m�i�� 5����C\��]f�%�F���b�z���O�����qq�RBF��n�ǋ̀i&�s�9S�'�zAA�z��-1Ⱥ����:4*Iv�-���$t�Ƅ�q���&4���*sy�W�1Bۓ8��Kxn�V7#A4ޝ'��nt�?�E�<h�`����n�h̬��	��\�F�xqĖ%+����,J������4��� 1��m�Q��S��l�M��F�+~�L�k����ϱ/���"�����$C.8����!CF]���~��0��y�Y:� ����|L�,=�⭕+W���
1�zv|�	�n������VӒ���%O�r���R���{֋L.�p�1�?Z0��p�9G�����p����q�<'���3���T�>��	:��=�7�J|W���/�_�g7�a_�<OIe�%�pnwF�8��OKO�,3Q���π��nx�|��3p���p��euS�%.��;����=�C����o�^gLKg��w���%.u��`�/����.b�����{�I	�;�޼^k�,U*hD

�rBr9:��Ī�"{���1aZOkCe%�r��'�� ^���������&쫿�⫠����nXEu��.�nan_��.�(m�TN|"��-'����շ�\0M\`P��_��C^�����_®Z� (|�1m�<d��9�i����+�bͿ6�kս-�C�
��Q�4��Z���d��MMe�����r��l��!-�`2m����N���;xbÓ<�e����u�(s�����5N�yݐ�1��:��z���G5����=4p��j!T�c�Q���S��~�uL�J�gR,,�Үa7y�C&SU�D��t�I����ҡSI��X��"��د���Ƕ�6c̋c} ���Ri#��T�����]�<T�"�u�}?f��m�����^�݊!�(׻�2/s�M���<{��T��+|��E�3���}�q)st�ޯ�6[ጚ�X�s�iW���N���lW�|$�g᲎��gٴ���y��Z������Ѝݴ��e3_m+n��Go��Q<�3'ն� ��T����ⷛ#����1��P�;^q`{��*����gg��[�<eCY�4sN��?�a��_�A!Z�h~\"Px�bR�S�/��(�x
��k�u��II"��=��J�X�H�uǑ��*+,�%�$$ҏ�����"�i��=]Eϯܛ�g}0��]���j.O��|�G-hnƖ���#×�3����԰����hܛb�@;�@A���Ӑ�rd#wzm�:V�r�z&[l*��zl��n��vmKa�v���[R�em
Y!eǮ����=6�(��|u�&�i]��{����g�s�+G�j��j���������/�ݏh�C�K�
��q���i�xܣ�K�[&�ᐇ�I�#��r->�ٿu��4{)����7�ʹ��JM��X��l�� ��_:vO	�Ϳ�ON{$�VX�BMH����g���w]<�q�ǯ�&]g��#;�ҕ�|@��h�ߣ��g������0��V��
��(�^��?-_��`�� �_�����K�e�6�9�R� Z�������<�!�
}k�u�r�����%�6N��&�ߗx�葹{�1�5�B�p�����Q���]{�D�V���"@��te+����>W(g"Z8���9����o�F��kU��j{�������_�($��rO2��a��=9Z�3��M��ё�&́R�Hh�#-*��E���q)�׀�B9<���<�Jӏ�$Q�-pe a����IV��#R�`��޳�� ����w ���P�i���M��>c��[��ߝu8l�������|[i|-p�[&d,��UeJN�P2Lph
�[pރY���w~e!M��H�)��\�6�u�a��D��L�dS�P��ZV��,�M���/o����\ǝ���ŪM����[Q�eľ���H���|pvì��V�3,)���ŷV^�$���Vʋ���4�l7=.Mƻ�^����wkK>0o�)�b?�2#Ė�ӈ?�%�B�NU�c\	��>N�8LU�ȕ�/_�n�3��@ot�Ml-�<���`W�
D.#��k�މ��#�W�D�ck7�$#�,���T��.e��[ NeR�����5����k/ӺY��4*���?��5CB9����vU������aQ�CE��9{.�R����e\?��Q��c�0�g���_�5�`c.�Ge8h���0�7�0������˖�)���=�c>h�k��Ξ�XedlL2a�M�թ��{�J1&u�Խ�p�8s�2>y\D��Q���Ϸ��X���4�P����������i�x���.<�L�j[����Jû�8iM����y2�h�:������O=�W��k<��w��!�%���B�e���� <��-�N�k_�QX���fv�T�4]����&�?qvύS��`v�7�����c+}�a���Gƣ� ��p)˂27��Z 3�����j��������'�DM��:/���%y��g�c�l:��vHӢy����c��x:c�h�x���9���ǣ�Ymh�*�K�e�F����Ei�����|����$s��agy�OuD�m��"����"c�u.*D,���6!�*rs!Y�
�ӷ�3��ȫ�����v���f���"(�V�c�1�'�])z;��8B��, r�p�{��u~ҳ�V)9f\�kf��P)+D	�zI��W��E���85;�J����6\9��a��,��*Ƿ#�r)����ލ�ش�Ϥ�f���7:
�1\l�t�&�d�~���g��Ri+i��a'՚$ U&#U��=NU^D��!OL�vu�<�wF�m�F�����*����_�;�P/�Twl�G���fro�r Y��[���X��[lI�?��	��`�7"�!Y���$��^wk;�-\k�e���	���ݢ�ʳx=O�1��k���s��V����Sԭ-��{",8h�I%m�@,E���g���\x<'��B~Ng֙��vZ�:�Ţ�Q�
F�P~����j�jZ*>AC�ףxX|�������g۩�]�����,'�6B/�Ư ��3		"-�e� \D�n1j�ҷ�iq����չ�Bͯ&?��H~;F��]�
!��;�hp�ƙ�X�fμ@������yf�� /�~�M��[�<��Ֆ=��7t�JK���f�w*#� ����t���e�	O<Tg���z��.�k�n������g:{��R�`@	��7��?���	���B>�-+s:�סrDj	6<OQK\v�FX�8��mP���><�9��ܐ
/�Ijڇ��-o���`���BΌ��t0pV��r�/�y*)BE%�P�_���C{��m��4���I�DgT�s
�QUw�s>�'p�M��)D�jf��W��k�A����_�7��f�b[&�-�pY�C��`����OҖ�}���=@����:�L�q`�_��,�%WuP�K�
6.�Z��6j�!7��Z�c��;������<8�ԃ�*��e����Ijz���f��O�l�Q&ާŜ3ZnkT��ևB���x��Ն�-��:�i�.;��	B��r�c_$�c@�ߡ��N�&mh��������5��MZ�@U6S�%��S�*�u�L���� f����;�>�V9�0OK���@W��%����G�>��8�� ���(��V��u�(XB���R+�y�:+5cZ��/,�׮P+M�I2���
��|����0����J��{{U�d�G���\�<X�f���|�j�Ͷ���0`7��ki��_p|�>�7E��Du�w�Pm�Y�"[�*{��eFɇ��Q7g�%�ṫZ[��M�X�.��;m���3%w�9�5��T��������%�-_X0��C}o�m��u��i�`@�d�+_h]d�Gry������tߍ���tB�>`��J��qa?�!�1��8D����Bm��*P�SR��s�V"��.�o�R�f�4��
�L#�죀���A��Orj ]?F�cO>~�.��k�l
\�G�k�ý�Iz:<�t��vI��^�����Ր�1���,O�w�o���1<k �dԫ����X�;�f&d).�tp�;Ǝ�"��CU[�!Sk$��ԛ�Rq[�{��M5�s~���k��<�e�X2\7����2E�����)�t{-�z�|��KH����Q���1w� ��u��яuʭ��Z2������<d�j�	{�{�F<Zk+,&�{x�{ӻ�"C�o�E�sc�`���͏b��Q���&�V7�
�m�p�~/ީC��`�sp�"`xN��w���z��^���/�_�ĭJ�oZ� ʛ���0Nn�g��E[E���=Z_�C 4N��D��f��,M9|��9�%����MK�L���x�$�b��R�K\��ݱ}�qB����k'�Ct@,�;F����+#B(��AY�P���g�?�X�k���si����3<���ϱ·�Äu���u�D���
&�f'��6��,i��u��V�����6_��[d0��F�-�Ctv������	���@��W��7]݆SrP�W d���g��">�qW
p�diY�tuɪ��:�|h7r�:}Rv�b�Ci�y����[�|��$܇�NO�νH��s��ly��ô*��#r2Zu
x����t'�b�=�^@���������h� y�h�{*��c.��m��r���^�c�Z�S��)��J?|����^�
�&D)E�G�b���U��~qp���D�rA(j���6:R��`
(�'���%E��n�$H{z�N�ʞ���Md�K�eK���N��k|N�d��`��uʸɫ�
��{g��[�������}+e��@X�����%��u�b��%\X�a�_~ժ����z�X�!��>��]�����Tg)���BB|aok�+]��o��)Q�JS<5P��7�η�HW�	���?�ϾpC�¬eyE��
@i$/��G,/���Hz5V⃣c���~p��9��7;��c�u�a��uH�f��n�,JL֟�1U�2��|�7�br5O+yCH�0�=ԉ�D���#sO����s��iEr�+�Ӳ�����v?QG�>c��]앁���G�}xKADAX�/պ�O'g�5�!v:�Dɳ����bv��n��3!�=��m/�z��Q=��آ (��T��.`O)���������p�0=a],���$!!I�3�Z���D��`�s�%��]f��迆Tp"s%��4�ń�g���X�*:�o7�R0�2y�}�AS��i�BVz�y�H@Eᐱ`��zT�r����d�g.mv�6�2����)�Bb��@�Q⩯{�LW�cA�f˻n�~Y6u��s��cbmC�\t�Z>ގ�@\�=�-6���~۶&b�fo3�j�[8�i���b��s�Q2
�)��@K�|��M?;�xst�iH���z4SHI�ܹa��dB�^\�34<��  V�ִ%���a��<^���h4�B|�)�#�Ų�m��V�j����$��{�(��������b \��Y/�8�%f�YO vD�V�8�U�������}D�/@y�[�u�'��X������h��؋O~S�O�����u�0�[��ȵ��۶�4.[�S�oK�F���r ��!:xq�*����P-Rr��w�8����0��d�,C"������OG�C����\4i!_ S�[����n�2��{N�}��S�.�d�����x4��<��$�	[��,���������~L.q֒|s26����*�IQ~��l�17|v _5�� 5�]��Ӡ|i�	�_��v)�|�5��x�Քo;���b����S��2�̇D{��ٴ���F]5�uǷ�Ì��rj��z��I�Ab�	>�+K3���D7��%���my�٦���'�f�9�H�����M�Y c�;#To˝6�B�e*$|"��tl3NC��[��{^H93���R@��Y@~�45k��$r��-���C�钺W�g�E�{ lK#�A;����;��XAZ�|��n��]oUǲm���q�����%t�	��܂{p����!x���������sjlz��twU�^k�9��wa;%��xpu@йF��oF�ft�7���6��������	i�?f��aLEz��< $~��S�&�)(�ӳ��h5^{C�Q����IKY*Ksۢ�D��1��t�m�c��/�Վ͆k���~g�����KQ�zs�I�Y�AX������%@��K���lf^;���N�Ԗ�ܘ��z�Q�( �Vp�C
q��hf%Ѱ�vB\ǩ7x�>���^�-��C�}]�n�;�9f���OAy�L���<�ku���<P_�s�}�yN_�T�o�.|�s�5U�Fa2�u`�4��B��w�Ko��t�����^&��1�K��Fʗ�r�y��,x�:�!5�-$�>Lz��aKkmi�5�W�*������~n���O�����)����6��n@)cU���o��6ѷ���<��Ktp/�� G��kx����_]��}�M2Q%/����"⅁�-�;��%�f]���̆S��$ �u�[AR����cO'p��E$�nԘ��ߙ��m�ug	g����B������-�k���=J�����ƭdo��L�?��;&Y�.��*[q{��;��.��M[:�Z�joQv���]�q�ș��6��3њA3��+jt\�ƈ���چ�rs�t~���K����N��B�H�		�[��������fȟG�=|)��}N�}��0ȗ��g��i�A���u���E6d���h���SD�p��ӎ���Q/�:��n�w��8M���+o����/�%��UĥN5�r3�=�l< s�~t���8f^�3�蔵�X3`�=�qyd�j�O�c��R�&'����Gg5�$�Z�Н	���������B���L?|���6��� �k7�t��n$ճ��E�N�4����}�[cc����"`T7��2����id�yv���V?������
%k�!�ɺ����Ŵ���g�&'�y	�Y3Li�6G�fQ�
���6��Uힴ�_��x�ԭj/(|�L��d��&z����l>�FG��|��.K��2Gb*i�c���\�'�T&3��|���r�`��@�'�p\V��B��h���P�0�R��)���E��B�G�����bRJ$��N`�p�w/g�KU��m�7�kB[:�_�>^��D��i��6B����1r3�+�`�*�D�]@Q@�gf]W.�BC\�u'���z���(J�]�����w�����1�N���d�dא%���춏����e8�f�(�N�WT���x��/�?=�2��
 ��rv�lA��h��#�q���E�qk����G�du?X�q<�f�ߝs�3��]	�������ImfS�w��m��y�F��\HS)6��.j�x��Vq\.,�Y��d���f5jP:d?	�7��L�(�Dh��ν��_��n����u0f��K�0��Ɋ��e��4�aA�
�Ã��s�CF�+Ź_��/-g����r��Qjd릡C���k�
��\�w�6�:�����k�u<�#b�����<Ϣ�Lf<_W�&es���;ښ��m�U�d���=�S����ӄ4�es�f����qb�nh�S�Um�M��y����4o�.h�֡>R���(�o��ENU���,�R0��4ù�#�?�Y���sa:�m�"c/4�:a���7 G�6�^D�)i[F|<zN_p�����AP�[֯�nܬ�`��.qg��\��"�������p`'�Vd�" 1Why|X	E�|��zv�^ə��v�cbZ(��)�
q��m��י��S��&�zVv-�p�}��QuϪcXE*�:�mc(C%"����aEo�CqG�t�&vӹ�_'k~鮿�>Ԏ�� ��<����JJ}�� ?Nc� ���P�����H�T��_�ڇ �e,�X��**Ƞ�*I�;^����Tš?«j�lWi��K:������{ǡ���V��Ҳ� d�6�&��~��\m��u������A<��2�L@�~J޿����r3c_��C�h���?����7@��RC���/T��U!�w:b�k�q�@9���[/�N��}"�HF]�I�u_Wg粕$�����{�ip�ܗ�:�\��fN6��~��bK��yd�רּ�Î��S�Պ��I���Ut����#3~��#�Q�����-ڶ�ԿN��y˳�/���$n���%���VM_=��b`���_��>G��>(�ur���jHY���f��F����A`Yo��t�b�	[ȃ�xu�s�N ~I�m���_�.f_eVKFdS��V�;Q�5�ޡQ��v��ˋ�����P���˙/��I��Pk��jia.���h"�#�9���=_���qJ�aw孓�h�Ri5hQz��eB��/V!Ա�`�EX�6k�#��iQ����Tc:G��̕�Wy����}}���ܶe��ٴ�U��<y��R�x(Y�ښ����Q,J�NT�X����nos�NE߿�ȂC�w+���H:4m�9���}�f��ڞ g��}�T�0�(5a!Q[�.��X]F�(�^�$��<�(���i̲~�^���cȅfy�}���e���!s�"���T��>�f�8re�{�����OsD�q��teTa����X1���ځ�(��q���wj!�dP����(��Cʜ�H��"l��ȅe�R�3�b���zEFd�}������9��5f���Y��Xٻ�����AK�4�^��?��Vc��\@����7L��ڏ��O۾fz��J��D'|y�{�	�S� :����,�#�z?�I�P�d�VxΔ�P�J�ck�3;#T ]�(t���
Q��G��&�6�������*�FaK�RNz#����;�L�9@4Z3��˲�M}j8�@J6;��7�MD&$��pC��0f��x�HW+��xX��Թ����Ğ�1����ۖ�%o[3Bڮƴ��H�����XO���X�izҿ�]J�dz3G��B�v���䌸)Ć�DG�ş��9�|>ϼ.	��2]�`����:��S���Z��*= @��~.P�g+��Az�k4=�t��Em� [⡷�j��
����^��
�����@V|*wc^���!���Ӯ�K���.��J�&�WS�]-��p���q���!S�x֋K��_>���Z�_�)��O�o�����m�__��8T��M���U�WG���N�H�@���-D�}��D� سe�Le+ʚ���Z-{���(-�L�҉��r�Hו8�E��V�	?��NH�L���#D�!��ƃ
 ?�u�C^'��e�W����+��>	�{��SdK����-���(>�4(�Cr6[FA�P���N��2��H����d?CO�h��'ϻ�( �g࿦۪-g��v�4GC1��=�\�������t�͊�+gK,8L�u���'m��S�n�~`��zࠗB���q�� ����ӻ�L�Ý�6�$�eOņ˃��`{�yn�[ OW�\*bky���"�NW�v��3b���c��I_Z�+%0��VQힽ^g�n�ܛ�h�3�^�jTrP�uȚy��I�?R�,C���������	����]�.8���5*��k��
O����YSK%�ߑ(2���QХ���}WW7������` [�1�:����N�|u+�ͳ��dڎLj��-��X�@m/M�p���sTD(vvƪYg���2n5{�C�����ֺ��u0.�֥�\��t9�:K_��>@d���@�V���R�IpT'�{u����!��_��*h���@��Q��`#&�C�I����( g����N�<9�%	�q
f�	��96Ͷ���eo�4
���,�y��هps#��BGE_Y-+�,ܠ��L��g:�,H�Tg�Bt��֊��w$))�׷Q^ͭ�����$���)�Q>�?a#��Nʩ��,T��1����aB�?�N	��N�W���/���~c"�c�HG:��x,Q� "y�W�e%Yp���C��'K���R&x��������S�i �A�+}��;[V�w�jO�@��'��	߲0[�<�|�ʼ��R�v��U��(�T��Hƅ�3�[��4��U9R�l�8*�ӷ.��e�����el8u�݀���i �l�����Х7���§S4��-�޹��	;���R�P���C�8Tq��N�T�L��[45��m	)R�1�������	��2¿��-**�NR[�Κ\�h@�2�:'nq�͖�$Ǌ�����LHX�ۃ!w����s]fR�f_���D�����f��Qc�##,����-2ۊN���l Н�+���#'9�"�׻U��BE��ڇ�e0#BZ���H�g7
���<�%v��mUc��8*QO*�B�iZf-�+�E�0�NE�҅��I��I��������7�N�Ɍ�/.��x�ۺ����� �H� =�I>��Y�����V����P���ɲ��o=W�]�h�a��n�vYĦKE������-VmH��.L�խ}�����u��?�+�7v� Uf�|�k
���|��)ۭ�D�X��x�W� �l��e&.P!��ᄔ�9qpw"eR�����Ĩ�H)�,��d(�+aX����+�
Zh��ep��5ͱ�<�C�g�{��?��,���K4���4����#�Fe0�|���C�H��h@����>rX�1��iZ6���4*�F�x&�IC"H��ޤ�zf�CCk�z��A��_5��Hm~ۍ�g"������%r�٘���y�k'����x�͜�|k��9I,�����p�P�S��5��D^���>��fǩ��Z,=�o���S�-=�$�Gָ��^x#a��r�������(Ԁc:��g7��I�@*�q���)��{��O'�@���n���!��4_㔯K�S��&���x���sėGsTw�/�2X
W��w]�j�4�Z%����8:���a�C��H@bvv�È���<Q�BC%�9:��0���:��@�X�j�A<K������+��hV����J�̓Yy����b��,e)a�r�ȂA`"dD���N�-�� M
�$	�!��l�,�kM��ӟ������e/��Nm!D�%���̈Ӵ��92�o$�@�}R8����"��)�`�� >������zHB�\�t��e��D>�؟���j��w>(f�1�UbE���̺���ߒh�%^�T��U���@>bm������)#)\�V0B��� ��EP~�ƱE�u��9W���w|�o�\�M]��Y���J]�s��E��Ų1�W�3T5�
�J�f����TT�1q~|w<�
�+��8m�m�b�ؐz����[�d�"x���� �e������$��
Ϙ�f\�F1Cc���^ʠ�:�OTG �z������P#x���o���	���Ֆ��\��5"n$�� ���X���w�§r_�]2����\f��(D�ޣ[�Pl	��>�3LԠUg������9�k刻e;XE��ZY
Z����H(u$���$t�r5��������ʝ
���/Bz5nԧ��+f���+�EJ;djv�)7,�|?�������	ha0kT�&����.g��&֩u{N��H������[�
�bŨ���I~�Q������])�ާ�1�Z��H�p�,�^�.��&���f���xύyA?.�?����f?���֯��}螽��pè��'�ϷhX�*�饠�����9J�
 �0|<p�,�tP [fS���! ��@F�'�#��y�P�1D�ж�����ΰ?��SL�����J���m�I "��o\�u�����u�~}mt�� �Õd��m���T��/��#��ɜ����kˣ���Qw'a��(HC��W,$�^���N�ܫ�Π�u�%v8����G�â��',�vr�h���@���VB�ԑ��=�ڗ܂���J;���7_.�_h�#/zÔp_;�0�m+]��@J��^ .�q�Ƀ��x�^�,�@:I��l4W�_������D2���=�\3���{�����f����Uݞa�I˵x���{o^=�����z|�
��g�>�-��9v���ȅ��胆�q��2��:i�����v�d�b!Te�^@AJH�� &d���5�I.;�9�sO�Ǫ�Z{��(T;��4Uek\?V���/V?����y���4�dT���-�@��n\����{l6B�o��*����5Wr�V�Y�Y7������į�5م�Ҳ:E�4b}_G{��:�����<��g����56?�Q�g����$,����].��rxS\W�#���M�V*8��l���m�&{�x�,5T�z~�b]�R��esMx��껧tG����DϞ~�&j�h�ce���'Dow�c�d�,�'})a{�&x�^�r��W��^ru�e/��M��v<>�������A�:���ܾ���傪�*�r�#��3�le1� �'�0�:�3�C����h�.��]��}��6E�i�֜(E�1��2��)A��I&y٣����w�=b��$��ސGMn:�#��׷tA>���3 �l?i���#�OIV�v�m7���9��[ejAx��7A��/���`ba��л����_�dp�>a�y�~��<�GkI����M��r?U��Θ���]�x���]�8��~e���(��|�r �ۉv��-�0�������b����5��^e�kR�!��Ν���(ч�転�VKP�<�v�Sw��6�?{Q��$ևg�\o�7�;\��N7��F;�T��B��ҌYl����=�Đ��/�C���7}O��/w�J�?�H���z�y N��q̴���K4>��q����|�ZH=ԑ���mć-��O������Y9Yz/FbT=f"!�3X�4�`��r��)��k�jL|�g����f����aIq���q��1��k�7w�'���J��|17��mnh�IZŮG?4�	��e�C������/�oh�
#�. �Ӻ�Y���t�B�ק�Ή�)���������N���zb�5���6���Ǡ{��A��*�Ζ�I���}Q٨<�)���a��$r��,�-��]�-(��A7���kɚ9v�1w��CL@E
���7�:�*��L#�[�u��G��<�j���^�R���H�����t�	%BRf�}�N%��
~#��lZ�'�4$i<�hp�-��a�õs84�Kjð�#%��3�q�4���*H��0)+:��=s���%,���N���MMq^<���w�8��$]h��tve%��-E�?(��8�NM�p0%�v���&�5v^Ϋ�_�K���{��sߣ^����r��r@���`FR��|Ta��QP
��!����Y A{�s?��������Q��S8�Ąf3̭�i,_k��h��ٴh��K�a�~��>]���چmm�1��5�/W�:��������o/��,��.�l�^g~@)���)Ȣ<�Wv�v��W����v����;�E�t�&V���$�6s����")���y��J�ՠH\��l	�2gng�����P�����Ķ��KZ�B�����G�F�6��'��&	+�b��8���������	<�|��~iw�8M�?CL�?=��,��P������%!��&?�Cv�_��fڐ_$X]HW��)S�-������1z��,��b�mx��S����gd"+�����l�$�5'GN{g�轻�@�=�����g(z<�O�'*vr��)���uS}��4���SC�K%,ˆ� �����
�.*��t�8����x�����~�e� ~H��ι�IV���HW]DWdE����|�޼1�"ZC��Z���	ot�g���6���`,��'cd���Z�������Cu�4(p�bp��w���Gc8��*�ܔv�m����i8���r��eVE܋\��@�z�8��`�6�N�����?��=�71��||���3�>�酄�|��$�xyFYw(��*�P�7�#��2��+%�:��/W�#�"�:��K�د�^+ʇ�"D~�E"_>�5@-wv6���[�Oi5D�%=����ܔS/��J� ��>�\/ۋ����>&>��Ν$k�B[������>���/4{��W{0�A���49�">ܢRCWc˅�F�={z��r��8�!
Y�e�T���ݹ ��ePZ���Ʉf`Fߞ�G�d���*Lk/+��W�.׵� i���x��+����l(�.g�3g������Jٛ��a*�pE���j�U©����\�
vn9�0�a~�yT�q��)��SS9s
��_�f2C�Z.��MN9ZW�ذ�n[��2���$�aX!��f2O�.��K����HQg��@WRh����?��E+}�/�Aa�fF<��滟�F8�����	��)�����lA_�A?[�>���U&!ͬZpg���8.��]�@<I��G��!����:F+K�~`�an���g��9���$�3�0!���r�L�"DI���X�_ޝ_ �̍�u-g*��������-��y���~7�'=R'j��#j��FE��D�^c�@��?զ����S�x��~�t軣r��A>v�V'��W�9�C�y�^:L�,�#���W��/ɨ� ������'�8�,y2M5!T���y�V���-�_�+�v̝L)ܮN	3�e��&@�t�Q������������Z��I���v/�c��K�Av\=휑 #G�G!���hҴ� Ou��n�A�&y��-�q�x�|��q��;35�r
&�,�~#*��*��i�Ő!��a���/�����u=o���ܿ<�y����|��]��:~E�˗��:��4���~)����Rw*VB"6~3,����Iy� ~J��V"��P��IiI��i���J}(��5�1�j�"�΋۵�P��˷B˂�i
�Rz�� �᤹>	�)�7��8�a���+�G�!1�R�[3�4��B��gӤ8�Z�����~JL⓽��7��y��*�j��F$�� �O�m6D�ŚB�%!T1?7�Hp�WG+�>|`Ql�����Jc4ش�W���Q���О�ae�M4��OD�Y�},g�;%f�*���W�sU~!�Z��x�Wg$�OP��!�n ���|�R�`���|�n����(�ٗ��`��4��	܄s�N�h:;��/�3�x������sH���"[b����o��%�
>,�����2�%7�4H��}��_����n�������q�F]r��y<0]�1���e���B�E�ACu�[��.�B叽�x����
�/T"+�[g#m���ȘM�0*����*i�TJT��V�F��"J��F{~\2�P�2<�^fp��1�w @�<e�0�|�w<�O���ߢ8LÓ��B<���UwW��)��P��є.�^
 ��jQNe�JV֚޹iE�tp�1��oV]���{/��[r
���Z�,<q�PP7�0�_���J7�9pe�Њ:�v�|���rkV*qY�+�C�tƘ�sTLy\g�������y+#�gD4� qy1|�����V�O8��%�0\���/s���B�����Oo�cF3ǁШz>�����ɾ\�1�|�a�P�>�@��լ$HY�l���}�r���:�R|U�c�x�l6=*�HW��M{"��@��)ڋf�m P��������w$�c��E7�x��[X��k=|��� b	���"C�}�<l2�q�p�����n�*\�v#�G��$��S�����=�{n�n�7Z��i{��f����uh�-�C�������id����1��*�Ã^*��Z������>R_��"��;����
'�m�1�����q;s��ʯ�[N1M/����~v}�v��Di	��Cpm&�F��e�=��"?����/�\�����Y����a����Q��k�;��7Ə�����]�/n�V�/�k��+�&h0^%��)ՀΕ�ц�H<z��)��<]p�rK�(�(�?�W9]Y��C]�ڹӭ���;�k�� X:!�e�K`�V��,��ѢV��i����k��A�`�h�T��"��O�v�ۀj����!�6�^S�V>��<a�����u�c�4�pR;憭Rak12Y����B��|k�X����?P�P�䃃Pny�Z)��Q9c&�yI�X�uǨ�B`���?�I [K���iBzI�	��'�
M������KaN,��53A��@����,�fo�Յ�s˧	��������6Uf^���	8��٤M�l��u��r݀u�4"���!�ˆ�ԁ�Za.�`�[A�����1Mϲ�*���XD�O�>qʘʙ�5́5.Z��J����I`z�"rR�P�N�,�F<������k�9��髣�I�Nޗ����1[.2��F yː�Bg<��KxI��n|�=m�`�A�T�^�
�QN�j�d!����?ZW�ȡ�rP��������P^�����5CԹ�z=7�չ~��2Xvؚ�U[r�7Dʐ���L�|pbֶ�Қ����YB0�X5d��.�p��vT;]MXo@�G̖�"�}��-��:I4�z�� �Fj-�@�23���P�
�&��G�B� =��e��;�Ӂ��4:y]���f�Z(�g����۹2�����R�8���	�
��H#�EG'n�+�z�n���>8K�����£A��$��C�)-ŵd{W48t)xʹ�T��N����V@�\8D��l6 am;p�e�]�a#��P�=�����.�{��xF�n1��}f�4˅��r�>�B�t�hA30-��*�����6�����w9��}
	��z��x���UD���c%�9�^�#�N*��=�-onݙ�x�Ң0��9�^�D��š/���"!A�Q��7��c5pϾ��I��?����d�d������q˖��>9��s+ڔ%�t09O�ꞹ8��U�q#�\�&����A�7P�ü2��Ӿ��?������t�5�| N�'(!��j�	C�X-�oW�<e��"��[O"��/�q� ���'b��N`V�C����ʟy=Ńn�e��m�>R�"��Y���^��t8$�j����^��m�/��&W�3q>&�N��E]�C&�=x&]�r�C���ם[�j$>}a��i!��سQ/�����D<se�>��!ˆ}�!��~�[3�b�_*q���r��;��g�� �j�|M���b�,5x��+��X��SV����3�OJ �y��'LDuT-#4����,@R)�~�� jkM�Y 
¦����/u�]�G�����_���y�rptv9ُl�Q��Y4�G̬ �a�ڀ��8��A�c'���4Ǹ�x�Y�l���0��"fc�
���'�B��cLg�a����F�9Ƣ6��S�av�-���@f���U��e���V0J��;Dח�&����KĬ즼�΄��{����[\�f�6��Q>�;��7'��(���Qэ��a���'5S�J�T�a �a�_��A�v��|<}��M1r��	�����:����� x_� �k��Lz~����s���T�eu��km�����CW��=�B�fw��}֦�P}_X����=�or۴j���� �=I��r��-F����M�\I�_����yL	2�)
�@rLܔ�5w1�� .o��	$���V��H��^?eN���[�:N��!�i��<ժ� �"yn���Wߤo�����wۦ����J�!Z���kka�B-�V֩�*���q(!6PZE��T92[��QZ�@���ۂ۰��01�:�+d5��Q��q:��,��1�<g	��&E՚;��n����b����+��R�Ckeb�`?�	�:�/D �*ԙ�q��~	@0 q�§߫�{#g���e�c��}���3Hp_�mFa��+���tx�֢P���`<',�.�̍K+r�c�b?���N����Og��\� 	���u����h`|����/!ړ����h��&��!�}����)͂�dm�Sr��>yg�<͟���qۅ�C�'_;q�YY��Q�Iu�g.C�(�-1R��\�� y۟�%?�U�"N��<�2g�z�NbQ5����N/�'όs��Ġ%UX-ʼ�Ka,4�Cb}(�~;?�%�?o�lU\26���Yz���}���-��!$��mb�D��y�u�T��ș��f��3sYN���+�:.�	q�Gǳp�T@��pM��*e�m�d�lS�!�H�}L�![i�|_.���Wb����/ux�g��]J���>���f�ƞH���r�q��Y,�y�7YauJ�����đ�,�3+3!�M�Q��#���0��=:H�6��yyx����tN̥�K9�Vp�6�ȕf�Kg�WIй�4��젠��.r.N����lP2����@�F�+��l �困�H-D�n�|%p���ԭ��( ��,N\�nB�;�.��ԭ��a3�P����~��|Q�0Nܬ�{1�g ǺC��n��1{�"�o����Y^���;�pTޔa9�5/�����A	��M�%+�&�dm��pc�)kTth'������u��ʌ�ϊ���BC)itk���)��kU@���7<ة(D�y���!@�Sk�_I�z�N����ft�-6�P%�������ձ޸���1��4:_j�F����KY�'d����7||�J>�}`��}�.�{���zbc²k��!�����եy�a<�[jPZ��gO��]BMB�ZޕN=�=#�ӳ�5N2�V�+0$m:Y�,�$���Qh������oOzzo��wA�+�lp��%��o`�7�_d;G/����!|�d(pB�����4��y?LU͙�#Ӗr�����Pr�*��7(��s���#0䓻�6a
�]2�g�I�0-KԾ�kJO�:̹3J��.��K�g3���ŇH��^��Rt̒{���4B7Nޥ�@,*�S+b^�&��o����kjDB���,���"�V��,28�c��Q3�p"�����|��9��y+>���BrY{[�_��lX�ʒHcr������H9��˓��s@M���ʓ�6ש�{_2���^S�_�ߛ���`f利�d��P�
Q
	� � ���I�1d#{�n�Q}�96e���A,����j�3X�U�����=#���5�ޫ��|�qw�AhB�J�/_�~��J蒡3�������zϋt`�}8��%c8`���ů�������l*,M��Y��$̞�(+��78�K:���v�5�m�An���k-8�6Ͼ�H�#l�v��Ϧb�y���"Ӧ�7W?oF�DK����-YIѳjk*�n`�l��%����ʆ�动s%e�$���$ �Т��N��"��gϊ|[�Rїò)h���3=&U�\}Ó���Q�,1�����r��r�M�B\4�P�"�A`8=�:E����W�F��7j�Ζ��;�ި���u��##R�@x�C�zN�;�,$r�t�*>���V��j�V=����^@�[;��뷾�K�,���F�[�Va���Y�m�N�����/����;7�Q#(y6���I@���j�<��K���2z1�eh��mE;+�6Hߢ��W�6�G��9:�˷�u�rWA��ڸ� t���mҨ.�=�7 �x�?���7��I=�M�>��k�YƮ�S*}�_*�c�N�)�y"$�]��M��7�u�ۅ<�؟XW>=�!�!�R��l��Uf�f��0��(#q2I�*<M�0�t0��P�@��X��=���M���������E�
�U�$������H��l����(�����������|L���ȉ,̷��8��*ٵ~e�Xsp2���G7�U�P5�1��6 ����;��<��z�\�+Pg�	1da�\�"K��ۙ���+�@a�7�%ع}]�(;��S��U7e�/�os�kGXz�$���\F��3I� a�*��X8���6�#c67�����=Є�'=Dxa�˭��q��6{��y�#��Y�=/k� ���N�����2� ;?��b	���;Ù2����~G!�����x�d�4p���X��t-����S\L��Y�8�HJG?d�4b�l�rl���k3SS���~RRif<I��@�Aj��>X���y�N*8��@�fF�0ĥ�>B�I�I"�5m��hծ�8̍��՗�1�t4��-�d��<3k�s*��~�X�"o;V$��
�>~�&:�F��U�hߥj���h���_��C����J�56c	�[/��C���"�R� �vj�����M���B1��ӎL��oR��E�B�7+D�4]�V�[s�_a^\jg
p��%��X֔���e���}c���=�-o��6���B���6����p�z��cZ�fv���?x� 0�Ә�F�u��麇��Ǣd^�sM��x��*��08����
!L�^xu_�9`>����KΌ��ރ���pv�l��[9E����&Â��]]�re
T�F���eT�]��֑��,�1np����&��pRP�Mk��B,(=��V�/V�T~��3d�-�Ȟ��Kp�����<�^Tn7)���YK,ǦS�N6uAii���4�@��-o��{l}e�RΨ�K��z*r�ǑX��2OXxM�[*n�O��e��+�W�( @���B�ѻ��\�)�� 4̷.\Y=�n ����u]2�	:��\�s?F<�f��2��:U<~ɒ�r�0�� h�՗e; u���_.�^&^���֑���$E�rp]����z>9���>ϑ/ �r�p~�,W�����\Y�z#���{|E���u���Xc��켻e����Jai)�S�5��7NQQ����aKš*lu5�����H�t����2{�ǟn�Do�lG��%|�Tp�����~E� �,QX��,��\r�/0���9k2q�c�7�b���6I��z�y����>;��Ϥ� �����p��R}Q���(�L{/ˆm��>�P :�¬�KL"@4Q���),�ϣ�RH4h�g�h[q��.��{�c��,s[��ek�	��v#s`���M��˻"��v�{V@��YvE�}�d��:$k'��������!e�;�2I	��t�[��L�N���%+�������WE����h��ރ�s�ǰ��E�U{���g��ĸl�W�1L�x�!���~0g&
��\"��ё3��y�����ZG������^9PR}B�j�>�����g�g�c�������&�,�����T2�F�2T��6 ����SWgp��)��ڷ\r�<O�0<��]ڋĥ�����~鵭%�x)5Y�E����N��l����4$�]~ݰ�BڹB��sk��0gpk�$ދ�q����U��(�?�Qr�f\��	G4�`��h$+��o�R�8�fe����+]�y_�t9��<(��+�هDH_N���~��Y�:̞�����V���<bq8�>��!�^��w�41� T�Xv"1�oE��Oۼzܼ��m����N�s�E����������D8ZҮ�~�����4_�1(3Zm5�5�TA�8YK��/P(��U��'=��u�a)��l�����w�{<��u6w�J�Lhr������P5u^1��U��ߝוF�q� �f@�5�`׌���9D��RY$��WI�٦0H��Ž����b��|�P:	$����ȅwSܒ�E��c��S� :}.&z�е�*��}�l/�ћ�/^�D�K�x���O�j�nu/L��o}���1-�D�ų�7��=�jasxr�^�ʞ��u���̉}����U��āi�WH����eQȏ��&�[%���4(Sh���Iz�Ǌ�h�2!�����)	��O�b��p�39l��������#�_S�����?����-��@5��Ĥ$�a��U��oV��ep��[W��~ ��Ȧ�,�n �+��-�E��:Rr/�ȼ@:I�.���b{�7ڶ����T�6�7j�O�J�*c����-���_�9����dT��-�ۃa(;�m�F�R��"j���.W3÷��_�=|WV��~�K�x����!9FG�4�ɻqo�&��m�#��ZpϸoD���틂WkO�z��φMD^��X["��.��y��=6.��h:�����w?�EFņb�1��;t0�@8�ʊ���ݽ���ȵn��Yz���QSY��5��+�����k;�2r&��4�-�jF�+7��hA�NA�<��8�%:�"�م$���Ͼߩ�G<J��Ȇ�����&&�D���&&�2��%D1�N}=z���e�O�p_��3Y���tٷ
v�↍���M|0uy��]l+D@5�no��X��OM*�+dx,�04�����"ɩv�`m����)��)�A}L�bX�A�i�V�5�2N-$���M_��Kg�,-(o -f��ϼ	�=-��N��8JŹ��w�;�}˼2y��w��,&�n)�}�pu�9A%��>`�wYBnv̡ESC�,9":j ����/d#��r�3$�/)C'����nbMz��jVÕ7�^��Ʀ�A��=M��m7 �y���78Zg}��������'>A4ʹ����2�,D6<��D,(���g����׮��9B�� fh���E)�d-��g����:p�'��t\���_�s�9p3z%,�Y�B1���Yc���<[��܃"}*:dT/�X85�#-���k��R^Z�ޠiKJ[	��x���$OT��6ę-ƥt����TNcdk�� ��U�ķ#V�R�$ƶ"q��&h�e�K��Z�[�WE����Z��������X��Y��$��FX�[Z�sIi��w�������;s���'ff�@�d�}]�_�c"J�ʔ�9
�.��B��;Rv�P��ֺ�s("�*��[��f"�P����J�=�Ӄ��ԏ���A�U�BX9�--b��E�x����7>-��^"�a����ӯ���D��Q�SB����Wp��䷿.���)�S$ЪH��-0�?#��j�')ؕP�ǳ�7m�k�7r�iG��;6�X,���i����� �z-��L��N��LnU+N�.V5�g���u}A��dne��EB\�����eN`��.;���Ɠ�<Z���XՆ�RǯH�Ar�
��qz�wh����!���Zprd&�[�g<%����.�˺�͑�ԗ��S��?�_�kX�"��rʛ��1�ݓ��$*���,,�m�P�������BtT �������O'�&pM�En~ÖU,``���6�-��=h�.�'��<�<��
��~����\�"v�WA�n�8�d��A	�uH��ĳ0�6�0s�A�f%`&E��.��X8͑
A��b+��{I1rK������緓DϿ��j��̀~3Kx�9Ƹ`Wr��*8��ೈt,a���;d?�R���Kx��-4׾q�(Z΂��'�Ï+�!�G�)O?�'t�!D�����[�.�
(�~O�,��"M�\�i؇��׭ ȫ������եG�!��e�B�4F+�D�>\aJx��Q/.�7]�G/���髺��IKݎ�{��4A-m?z�I����	�bE!����(1?�,Zl$)c�)#�)���n"
Z���`B����q̷zS�y�=��[��vC�d�v�d2!�����w1�4���}�	��mgU-���J����E��&]�{563f���������9oA]�9���C���mϳuw��G�W&�꾊
��5/�H��ٿ}�F�6B�3����hm�ݏ�������J0��Ϳ+��fTr��ڦ������{�����^q����L�n[1�&��8� R���tz��2Z�Ē���%+�k
�d�F/	y���ۅ��(K+�M��Tm�;�2D���Т�s�ђ����p�V\G����*�1ٰ�����B��_~�Jс��=��?��d� kV}�cv+b�u8Ֆm.��CqY�(_sp���=�UW���ͦ��H!v���Mf��ޥ4�xz
��ӿx�Xt��!g��G��sT�e����'��Q���$&
�R?q�բ%�g���Q�Je���<.gc��cvAI�W�Ap[.<T��	�lZp��f���T@,�cr7u�Z�#�P"��@V;�<ߖ��԰p8i��,Զ���s ���طQcW���x�0�*b�~���Я��8gc�Pfe�Ζ&c'��(u�|����Җ�2sssט��������:#X��gIKڮ�RG1���Ә��$�~k���Es�x"�l��0?���DH;]�__I�)ݫ���{��?�}� 
��ݢ�s�Fs�f�`|(�+*�r8>�2\/��1�;���.uU��w��źwl��)$6����x�EG9\Z߻���	d�	B�6v�:��K&�[���'�h��;��5�濾}.�&o���L65�A/�H��S��� ��K������ԍ�TG���$*&*����?Ê؀�efg#!�䪣DȢD�<;�L�����(��Ԯ���[�� H��'�{�3b�0�����K��}��חl$rl$�z�~
P'$�`��6¬���MF�d&�D�T���
��v/��?NR��̋��hv_���RT�e:}R��fNSVUS�b�VQV�������T��l9���^m7��׻/ο�t����~�8D�<�Hg$����˩�"Þqn|��q|6>P�P�]q{k�qw���%M�%-+[��8hj�����]��Y�޼h�k�e} 2|Ib�u2�;�����D���E��NΝ1�;�
n�������i�rR���̋����J����-�|r�]j��BMӚ��O�99rH�J�N�GG����''m2��(M��C��P�`��Ay��"~���6Aά��}�ee4 ��x]���3����-^�d���Nd�jTb���D>9HJ�4Fj�S��V����dZ/�?��L�nngƱ�����e�����ҁ�}~�pe�?�/Cj�k_	��%<�V퉉��pB�Z$>���͜����_[S���N�W}ˉܺ���SFw6�@�n�ꃧ?V�L߂��EA#�(Z$g���
C���I>�]c��Ô�*���r�g��9Q�} ��^�i�'>���	ݺ��A�w�����v�h%���.F��������͍H��i���uLQ��H�I����-���9U�	��Pi"�TK!�PR���/�~\t���q��pkGS7l����X"x.�<-����v���V�;T}m%*ZZE^r�4�����76�>R�ϡ�f�T�(\�����e���|	7����9,�G*]1�Oq��1��
_
�ڋ������ wYX[� vz�h��>��1X3����i�p3�E3��
���%'Y���^��_�w��|bbq��Z~�����,�W~(�o����
C1��p�����:���V��b484���2����?i��ڴ&�;IH|(���l�x]h,��,XM��yT[�f/'��\(`/t�P^�t?+���.bB/($��ʪo/��<�|��������T��N��r����{���O�
e�@G���r� #�_rd ��b䖰���݆�n֭8t�^�*<RQ�ڿ��Sa!b��V����`�sd�`!�N�Ô~�ԡ�|-e����=��3��`C����ͬ���Y�| �%�U�I
�U���
������2���lq1
����`߉�>�5>���\d�ǝ�k~r::���^9%%�l���I��L;�35�(_���u����Ak�z9K��]s���X�P��;�-ҿrt��B�Ś�Z�0��w�F2Ƕ�/�����l�p�T ?�I&,f�������}����Ѕ�J
�g�+�D��a��$�f�Y��˫����K���&��nkI��../�T'B�s�R�m�æ��>����館$�Z�E�+ZOg����~EEE�A�*/�����x�Ӌ��7�Ն�1T.Ԡ�����-fht�s20�|!���"�t� Hy��Ϲ�B[sv�H�{z�@��A�<���L��2�)�.����?h��K-b�n|�^ ���0n̟����v�20�m#���s2r@"S����i[��a���l"�mm�S?��ɵ:!#��|7����\-�la��^.$$Do����ӧO�xџ,��T�I����
�R/m���xyC��LꜬ�).��,��qhhh��VH�~:��H�����Q�_������-��E�������Zr]��|-"mr��ŝ"M_�k�~P��Pƺ�l�FCC۹~��!r2�v��O��5�:�����ɰ���n��lM������}���H�cJyyy��^Q��x
On{�dS��g��竬��%	95�Gi�j"0P�{AЉ����+��3]�����Z$8����-Z���,--��:꛴e��ަ}:���N\��>����J�+���n������fc��	�,a�A�˷!f_�"_S����Vß��n�7Hѭ�W� h���s���:���VeWt��P���:s�8��8�/C""Я���jfY����[�<�JKY���pt�ZYY9Ǧ�i���3�V�JJa���0����|#�/�US����~���*{�Y�(��wrRc��-�Zm��A��砾F�p���P�ԓg����xl�'^����R�X�RbL�~:�����%,ꡲh1�{��-��ay�j�3P^Pw��ܻf��O3R�v��L��k>j�.[�+��5��c5�fD0"wDr�����#��� 2@Yzz����~���
�>��|2�u䑨��geIPM>$D�h��G��VCI�uu�@��ڎ��&���_���"9k�G�]�?�V�����+%L|�v��ǌ�chln�Z�j���?"<U���=�V��M��on�~l��K��1_kQ� ���~ϫa,0�
H0[�����'�˯�"))	p���@cX��9l�g}��?��-c�iD[s�O�����Qr�@��@&RẬ�{B�?2���k�5��4��ɂ����WTPS�?;;�f��#0Ͽ���D��a1��������.,�J჉P�_-;�9�m!j��o0ʭH;�2�Ɵ~9���G��<ݳE2�Y�����gg?HSt�Kb,����3���V��x�]���l5��3��>�
��^]�8/���w �A�-������I.F�ɬ�!Q.�����k/�<���zM�����/�u�6��G Z>m���=��mo_V^����+uN���E�.�gPI4_��˧R^�#WY���B牌��^p�4�_�g�
I0�!FŢ�����XV�4�	�(�nU����FD�gi� �5:�{���������\�';���tF��N�;@h@@ N,��,/ L �81�ާb�F���7����Y���x�'WWW��[�M�� ~_X0�KS��Ÿ�|#N{��ʗ;C�͍����.� A�(`��2lzj��;�y��]J+���? ��U�W΀y �<��k�쾀5�L���e1V�wK3	�
�	j�z��{��;�ún�ݞ`C��/�&9������{Xge����g���� �_��9��,��d�ǀ�Y�s�҃z�]���6���{���:��_&m�C|�e��>��p9�
�p� `r`�&&&P᠅��YT��������M�x�Y"��,�ul<��w^w�Pd/wj�jo��!�E1�Vt�&�U���҅PX�1�8�%Y�F<����J]PE��~h��!e�����=�|rc�������z-M���>[q�~�ſ�#u��R�� ���c ##C��y���@���8�gP|ĀM�HY%����U��([�� ɪ�1��<C)�e�z�r�~t��/+��ʊ�ߓ!$8@YTBPd)�efH�S��y�����JT�g��p 9���5�{'{rm�H�hx,d�O�z"q������$��>a�@�#�Ⴠ�<�@��J��*?�!Q��,��d�ŋa(��r~��8��Ǉl(�N8��+m����ϕ��?VN�
m�R���wH���ߜ��Ϛ3���R|�F`��h&[uO[Y:��H��v}��\��=���9@n|AB��P�60��;�A52���82��7�N@�-ԃ�-S�p��L%L��J-�\�u�N[kb~>���vr}��d�Eu��	�	3����(,d���ZΠ�S�<��F�{�r��.�����n�sw�w�`�
hy�����4@1�e��M�FH�/�F�b��??\^�BgG��x�=�t��w ��GF��h��-#9���|y�\���dgl�,tB��]����1p�6�nP��-e��-���C�Y4�;@s���hq���,/|�E)�����/EZ�zzd�A3��*�|���|�	����e ���Q�<6��S�۽�m�}^价��A>)�$ ���C��gҴF|LU9�#�&@���"޿��N����g%0�e��.�|��=!= �|j����T�lB7�.	��=���$�F���v�l����e��WH����_�=mmO-��L^jh$�|�}zx1H�_:�@-���t��Hmvji)>6��� .u�ȃ�`+�o?~��?�]Pqr"4��R7nc�j��XbV.�9o||+?��Z>cKs�Q9���q�q�-Q�k�uQj��Õ|_�$�h� S��Dn؟L��ᤷ�ف2�,�l�rά��'�{
�[C.�h�	T��)���d �5�����K�,!�`�OЅ
��a��o�w�X1��L}0��G���>PWE(O�C�����1�1��U��~�r�����y���:L��jB���h�4|^L>�������[�Ȕ��}E������A�v�fo��~���^#1(--���DDI%����$�ÉEvM�ȑ]�+++S���)bSY��F�-P� ��O��s)N5�$ �g�Y�
#S���WU �$����a�5iuՔ�S��k@O����_[��}}���<���p:��r�?���4�[��85������u,�5�}`� 2��5�<p��0|�,�]v�`�588��<ؾ"�SP�u�.}�҄���B$�>Ed��
�W;Sz�.��יcG�?������%�|>�e�U��]���(�+)�ZM�}3���v�)~���j��Z�8�&r�W'k�!��'WsД?�\��ۼ�i������[^�6=*
�;^z,$�i}%��_j9�k�����&�nc���~`b���<��OAH��}1ߜ�h[��oUke�ճ�f�����h+_�l��W?���a\T�|�Թ^	����a�����K�*B\�fH��a�G�98 ��q�TTT�/ᴊ�C}��%_�Т�!uG*�������J������L@����ݒ�E���L�y����A�*+KK}��?��,G3��L���۵��|�A噁�]HJu�,t~ 7�Ȑ��jG�(i��w�����+;�fՀz��6�ݹ����o����q�KT\|�\��31��^-j�rn���a0��M3�������0��GK2Kj33T겤��&�wt4.����V��4I$����:)>1�A��>�N�O]A����]�uq*���\������c��Q���zƶ�~3|�R�y�AFF����MKA!9��u�i���b���@�e)QQ�u�C�k"��S$�>��,����<p��x���¢�aO�J��y��"�I"A\�a�� ^����H���М��gܚ�;z�s�M�8鎈.闚���i������L{��?1x3kU�hS0lqp�8����a��{�VG�!k]���{�H�V*h��臣r,68uW-�����n���8 �����k�%'3�_cAja��7�������Ff�{%��F>������-�7E�h%��.T����Q��S8�q���G$�F}�>���0������C��n��-�kO�v�ѧ���e4�(22Jb�򓝴�M����ۚ��*%r��C�׀���M�l��р�mT4�GDKr��J����T���������@b����\>t&/��YX�-�xfff�_�/s��Cn��'�y�0�ߔЎ���$��Hj�����GBt&��)��<C(������y��%��i�e]�얚��fk�~}6��Vj�����M3���3�����G��dxN�b��S3��Z�{����gai)��N�V^U��̞������M���Sh�H����)�&W\�j��;
���燇[���c�����g n\�଒�ڃ�Hn� �h���[��w��٥�,S��z�,V]�r��f����F��(tK0ۆEֶ���E��dv�(�r\&D����g>N'��)�a�]cc��z�$����'�P+�%a�F�d��A��gK�F���.����bdd��x���,���n�lr1�ǒzXn��+������(���T����>9��!��u��.>�eKS��'	��9�D�������g�ޘ������
y���ˉ�ω��Lvz/�J�V��?�����kSc�;�m�������D��`�ɮ/�dH!3y�����핃�8������M9K�J��9vTx:�1���N�s�
˟����?��^��H���*?&	��R
����|�+Udh��o�x��y���T��nX&2��1Tύ�>�W��jW��p��3"�^$��`�oɱL�M�u6� NF-5%no��j�4,��x=�+��, IJ�S�U�mӰM�,w�q���a�k)�N޽;�H=7����Ǘ�9oL�9�����%�v@1Vӽ�[�A��Y�6~������e �{�]�_k?`� ��zs��K���|�8;�jkN�A+��.p��$�^�D|���u�{���z����uNZ˛��4��:�X�Z«����ӪD�5S�Hӹ�0����iZ�����Τ�
�zA�����8.L*4o쇣��5�W\����͟�(��ĩ���N "�g6%�@<I���g5�A�%�wof�K��P�f���3�/�l�<Exo3ݸC�㕃$X�շ���I����G�~Qړ-q�E"�������� s�Ȫ�=�#����d�]�������v��Gvo�� ֯ud8��_3,�k��ʛ���(=??/#��HO@o��]�y��x�("#����2�Bg𪡣#�Y(~��Q�����`�B���A�h��p5V`$���Di�z�z����K���6�s:#m��T4��tC������ٚ���3�B��殫E�<
i�7{�f����_�#��T�
H\/{c��zl���ău?�UѲ� �+�����Q��1Gٹ�H����K��	q*�vqI���oi�5�~���;MH١S2.8�.}^�V7��'
5'G[�>'$5����~qg�`F�mh� |J���IKmxق�,��ڪH^��@H��Q� N䑤!�T��}}�$c"�e�UMΘ@Xh�@G�o��?8F��ߍ0/d{�G=Np*pM_\Y�\�����6������i�T��e��/>�]o��w�C%..^�vWO�_1w���#��p~y�k�V�9]oj@W���36��P���/�^��<��*ډ��?6=S��9��b�р����.��n�ܝH��e)�/�]�F�FZ�?�L9��F��� k%}���~�Zjv#� ���E���Aa���z�-�my�5>1�=���wfyr�+%�$B�~��6�C; ������R[��[Dp����sÿ�����|Qro�iZ�D�ШvR$)��
l��}��T��?~;C��`��m	c�۪G�?]�%E�
�	�R�|�8��¸�,�0*�b�������`ڌ���dy-��o��"͗9��j3h���b6�&�*Z'}�P1�Rf[����#c�dZ��oٔ��[�������Xl��c1�r*��?��d��_�>������ bK��Ls��:��#��e�=;���$;8�GUX/uRi��8�B��:N� ����)�;�W��!K�o߾HPp}
��%Y�=��ټ�3�����5X�����&�ɟ?��E����|��#S����XA��үd⚖�_�o�}�����S=p�9��ӱ�<C�!�����(׳{�oZ&����N�d�]�[��<}\��������<X]-��(�����K�"L���Z  C�]Y����֖��v���������?�(9��|����1�q��ce��,Dt�J�!m$���O�����r��H�V���J�W�0���B}�������^�Vo�P ��x�S�y�eQm⯂d�Ν���ΛZ> ����)	u�ժט\�&=pC-�Y��y(���n��3OcRx9�����k�L����� ����d0|@�c���E�a�� �x
䄊��Vc�q��������.��ه	��B;��u--�KM�*,k��v��a���(o�(�zP�=���c�E#��� B�� �m�X�q� �b�o�Y��%ź����8X�lv�`��`�����boT(Rf:D��cs}�-�A�������4M� �*�K�F�x�t:� .���<ý��Qj����]�0�����q�̭h�����p��V�c�/)$���*��`>jM%֩�g�l'L2��lQ��%�0�MK_��u)�R��tXQ�Tua���	������Ĺ�z�XG <�����@[�*B��&w�J����)���
tӻ��'K��f�!��K�J��r#���4����?hN���W�I�gw���XZZ]_�O��x�vO:4sDs�'��5���-�������nc�F�t
5O�u�����,W��"]�ۢy���J
K��*�
�����9��U�&���'ێ}VV��jb����QhZ�V%�7��b\�
A���r�TIǖ1V��,9�O,�&�� q2�\���p��a��E�\3�3��s���D����ؿ٥��it�GGH�_�~)�yf<��0$8r�ӑ�/>{!ui�%�K��*��Mg�~��|~�y�$EZK��]$v./}���D�<�(7�㺎�Ɔ$x�CK�ŋ�&%�Oo<��bE��Ԟ�!�@�w��:�bP������C�Ie��JYtߣ�C��z	��1���%�a���+D6s��7�`�?k9�[�_�x#�Ǹ���%�ۧ-Q�^�~USs���dv�wc�8�m s96��B��b���*��`�H4��U�� y��"�jZ|}s9��u̼/0���XHh��0Y��'\x����KqB��g�"'��J	����=�T�_�i�f�T45`��������K�%2r�m��w�\��{/��d��yf�6���̺����r�=u�6���،�t�5�m��ᐴ���&მ�Mj�Q��r7�ߛ�0�I�a�󡨙�^�ͥw��6ߓ;��m������&/��o�P�nu�~Pf#��9�~[�������\�'�iA�W�S��?/��, 
�c�wZ�u)Ƙ�1 �c�\̬����᎔)���N��`MA�9�~	�*�#�����H�� T~��y��*1(icH䞝;tbN^��Gf��z���o��f�>�$���nK�=�r)X�ݽly�nD6�P������&�W%�O�!�������42N۾VK�c��fP��9�菱��� V��2ݜ�[R�f����@�Ϲ���S���؜��S��Ό&s����$�.�,4:?L�t@C�?�������Cd�R�vV'�'�L��%*
5��")�x?��:�z�GJHMO���-11�d���@5�	���.L� c��^ԪK���q��g�T���v���!���Hl��n�~�����A�> ��B}���%�uV@�eu��s�"@z��B̅��Ҳ��s#Ѓ�ٶ�ñ~��3�z�f��U�O@ʮ_���j7�H0�{f/�ך�ĭHj�Ό&�q�x�W�����
F������d��N�7o ��%��+i����Ǭ����*j\��H��|?v��W���>?<5��X����\�%f��B�����˜�!�;�cf^��]D�A4����X8�I�H�XI�5�<���ur�{j�@@-�e	#����zp�т����:b�c���ZK�o������~n�D(��銵�#��Ś�G��P�.AI��'���z�:2����f-���BF	3�=U���&�5���AT�e��H�I�`���%���l'��y>W �[���#ꢒײZ⏞'�m�B�3Kc���T�R"�����I�>R�m���� �wn��f3A,�>��fo��~3�dV���7�ڌac��&k���kq�XJcZgfb�̏hǁ��3���^��<7Y�9M9�������[�%�f^��?�Nb�)Z<���fa�MZ^xc%=Q��U���{�d�)8�ud�RJUu�XX�W�����F
H�܍?�t�
O�&����+��b��;���~[jM�m�x��	
�;�b ���i
�$��S#�{y&��5`<��I	��!*�E��0�)Q+M���p����f�4���0�1O*ӯ-�����j C�h.��+fC��^6 ]�&9�5ؕ��w�{g�Xnnj�ȋ宬�~�^�Ѵ�Q�\��I��|l��궡�}y.DC���SԚ?+����%u���[��s(���_t2u�m䦒���
���"�Jd3��xo��mR|���\��%��,02k_�K/�����gQ�,��b`�i8Zyi�|��7��YR�f��4/i%�Wm�7Q�1��l]�&����@����=<�tq�W_��F�V'Z��[�Ɠ)��%���)��n7��!A��L�Y���|��V��zr��Э�%u2�o�46�>T��l�'`2��m�����rFÛ�P��GÅ�"ć��a"��$��"���Y���c�[��Y칭�TtlR�{���]}8�"^����f�qer��B����:��Zn���-Pm����@<��T�����AGs`I�8,�A ���-\҃�i�����a�C:����+��2w%�A�,��ky��}8>�$]]]�K�"�7[�O��ONt��-+PF��ѓ��9��ܜ%u�Y�W�;�8rGqt�a�E��H8O�ͩ�n�΀���`�M� X#](������q~̑2z��"D(Y� M@���۞E#|�Z;�x��r����r?d��	x�I��p��m�Q�?<y���T�4�P��|����c�gk�7��͍�t;A�?��������ߝz���וF���f������*�
�9�XRD@����7��꺫~3�J�kX[�
���7S��U���f���r��u6�K��N�u��^+V��旷n\bl���5�����e�rP�&��o'c�#
2����4yR��d���A9�ڞ�2���f�G�1���_��=��P�"}�^!D��A��&�����nΪ+�T&�44�m��=Ɂ�}V�;�B��ν�[��O�[�s@�wO�+6�@Ec�׋��؎�F/uF�D��'�>���:�ލ��f���:Z���6��������ݷ��F�	lف�Z��v#4�ΎD})h�J�:�[�o�#�$Q�"2����=z���&8ۤ�]��:tv AUuڡ�@D�ֻ����	�:�K����f�ic཈�(]�@'���4
Z?��+��I.��Ӆ��ϕ⶟��>N?y9
A�yN�ew��1� u�b&������\D8�Й���������đeҐ�.Ӓ�Upgv�І;�=1Qe%R/b���b�z�����i]ƙ���N�@�����H������&,k�]�����b$��쿍�4���@�^��M��(8�@���Y��6eU�*s����?!1���1֜�l�W�U� 5���Vi�Jι--~d]�.�%2���>s�@3��v������^��٤�n��]��7|C6F��>����lkz�g�v3u�u���[z��2�3XM�6�Ѭ�Cnޅ-`��������x
�������1��נ��hf*�;>�:W�wT����g�[;F����ޤo�=�2��W���kŭ1��/Ɍ��SCG�~��[P�A=d�HQ�v�a۷������IO/ʂ�W�s�IK.������5Y"�'/�B��͛��U���&�	0n�׏����r���l�:_��\D�w�<��� =�^	G���:�G=.���`O>X�#�qC��yl�A�a��*��O�����H=�ۇ�j��z��	uӍ���}���vZ��x2���	 ��S��n�p^�a���N��O�4�9f=G[��a5!p"���|`���y�'J��a#��~���(��p��F��������Z�^�uE����*��Ɯ���Տ@z������"	*%r��O� ���@	*C C��0~A��o3���υ��a�����"]0f��i[����H�@��������\[�?�ILld��C��X�3u�X|D�)U`�@�{uI�.'��ޟR�bE�e�R��z{��߄�t��S��j��o��RbԘ���B��Uo'�Q��� $��˧?���[�~���Ii�%O�@�P~�e?32N�|3	��| �*E�{h��ɀ�x���ah'9$�JΈ�j� �������~K�����Z�Q'��:��Q�C7q�k���US�@J�����w��lT}�)*�"���	)���N���`��t���j�������� u'0d�s��dl˸�:�.���޾�/����5r���f/����}��E���_6aV�Q6�?gd��l�ߞk�1Z �	s�CP
�bSb&�vڎe�����!ʝ�'�q�s����m�)}��@��r�ٯ�G�/���S>	�>�C4;�k@���p� ��1(��l���l8{qQ� ���[k�#�P[Ǫ���ca/k�k녛�]�<FL��Z�31�-u�7�d)Kg$��`��-"x�7��52 �w��`эȡoM���L5���d�H&vJjD×st�K&���t6K����]��+{�Z1<`$
9�Ǻ
���`)�����-;7`�ˣ��C6Xec++���py�C�����|{�M��uܥ�t�O�Sb���w��>{�L�w�E� �H>a
�	 	��ۤ�Z���;��wV\�;Ko+�O�m�޻���7Y�*0�ك���%� 1(tE�-�]Aғ�;����J�t�<E �d�m�_�'!�=��m���t�׊%���iJ3�+}b��Θ��V%h�_�*H���ئz���#��@�=E�D�3�9n�l�<��?b=#�N�E~I��q�J�>3�Ybs���~�sh*��-# m���x���3�,ٮY��a�İN݊s?�����V]+�h�+b��w�V�LepKg�ڵm0��Dx�"�BаT�˼��pt\�`=��k�� 0��O�.�����#��Q�����}a����xB*�O�{���q�R��]� M��0V_��ӽ�R����,v�� Vt��.X+&^�b�hI���4щц6, �U|k5S��*a%�xIR�b�����Ӵ���y�HS��%2 ���r�Cd��/ҦbZ�e�T�3�d�"/^I�w��(�w�A6vU_t���$b���!��+b�cn-����"rD�½Ď�ϡ���&e�i�B��4TH�7�y��(�??�ƜI��b��2�KW��S$�o�b�� O��,��5-QJF���������w���O.�ļ������ �:�k�~zʻA�1�*���u�8��E��r�� �a��ɦдJv6�Q�����Z-�Q4�9\w|�!�Zl$��q+.��ǁ)�f�X^h����`i��!W�Pmx�z����=�-��KjDg����TU�(��o~����_%���%=�[��~�ԩq�� ͳ��h�����5��mb�.�d�������x��Ԡ�\Z}�IВ6������]�(�z,	��	ʿ.N���%�����o�5o�2�+y����ut����.��{}�xҡ����>����/Z��p�3���̭�#���qﶎ����q���G�K���2�{C+do���v��� ]�D�	��`FB�]zr**&E��L$�^�eWS����m^���SA7na���<����p<j|�5��R��{��F��*p ڡ\�{\���V�%��Pγ*�F���4^!!����Y8L>?Js�fm�ds�����0��b^.�ժ�q�+I_<=��N�����O��ַ� Y�rv��&#��@[]}��+=��zt��Z���z�#�Аa*?�	��|IB^j�W��φ��bJݤ�d�C����R�c8~89�$��H�P��_����P���G@U]�R���c�!VS]#/��=9��e��E���R�s�E��i��ddd(�<�RE�|�-��yWqr������ZL��T0�ŀ%��0p�I�v�����&##�y���\�T���|LB�ʭ���	���u9XGG�)�a_ش��D���"AWF����h��6�!ċ�Y��GE��N����]��Hi�����xo"W^^~~uUjž��!;R�Y��WDk���$ul���%�'g
�U��R��K�t����.��n�*KDb"�@�Z��=��ն�
��������_<i#�@�9~]ܠ;�'��Ĩ9Mm���a���! ��r������Q�����'�V�A���<�f^N�U���c5D��a�r���y�_o�y���Z����HV�Ϗ�a�#�|{�k�~,�jD����5l���%B6�4V�B �q���dzu^
��q��vrC�U_ׯ�1�y�"zz4qr�{�jyHn�;2����a�����e��<����A�E�g�#K�a�r\!b����2-ƥF��@�L+=E�iz�J�%�T߫����TVn݃�����ܔK���4�/�����h����{�X�D�gt�h�uZ��44�7�vefg3�h`�"5B#��I`��O�����p��|��0�B�$�$�Q�<�i����DJ��d4i�KHLL�(��M�Yv]x^^�DUMm�'���*>5��7f��͢QI���

F�_��rͳB���W��!u7�$b�l�$���v��W.٨�JB9`N���.����)�P,d���=�'���%��?>Zޯ�{E��<�w)c�>��U%���	�&�V%5Z��H���������گ4�n��ANN:c�C�4�'x��i{�g�f��c��ĂoO���e��9�w̻
P򾃣�ζ����>y�B�����4~QQ���#�����^I��y�=?O������D0����:��0���j�ƻ�`�aB� A�r0r��$�(�0�ak�#�[��Mj㏇a���	����B~Z3Y�}����_��,�Q�Y����H�\y�ĻM�/ޫm%��b��ts^��j������g���(yJ�ì�I�x��.�{����0�b<ebN�=�4�V�Z��`�"R��70c*��$���R%C/�Z���Rš��!�߃�����㹫��_���x_,~��%���8�N��P��&�<�%� �3HP�o ���T�uTT��>L���4H	H7"%���]HJw7"1�� �Hw��]������uX���g�;���������dA��+Ex���&�g.�_Q,s���|w}�E"/���5��%u �6�2A�Y�����[.��V�ݫ�Ӌ��8!%%pt���POMc��H�)2�W�������Zi����E�$T���_��2�d�(��	J�"*ŗ[�����x����<E������¤�Γ$P_����` Td%�9Ax!i����>$���<'�R��/�K�Q-��$'��3�z�����s
���<f���Mk���x���ߪ�_rqPl�
l��F���y\F48�t*i�yXn{�>���S)-Em�sZ��x6+A�fk��jGl���`�-n�����h�k�t� �}*[lq��N�).��4�?+���珽4���F�O����i3�}����bG(a�_]	�M��A�J?rmI�%T�̖0�#��Pa!��|!1k"�Te`}��)7<D93x�Ӿ4����x��oMt5�v�ޑ����l�H�0�P�ku-��H|��вQ�:{u����W�����]�����L����Q�I�Z��gh�d�7�#�J$sss��������n{9��p�f	6z�o�Yl�����<�)��5l����^1���ؐ�۲*w)]T�����JY%l�n�l�3 ��ǀոG�'E7`��C�T��ƆϮ2Sͣ�> I��'U�I�D9 ����h��o>ha���!E����v��1�8ٔz��֓�ϱ(N?��#럥�1 �*U�{Q� ����c���gu�Üb���%S �pt\�E@@&xam�������U:ј��#L���ϕ�F���<پ����k4�%kD�d�t��������HZ���8C��/W�	��z�(:�fbb"�!~ˏj���Uh+=�hIl�7?O�Xl��s�ʟ��8�Z;B�_F �q_'����S�
���
�����̳I���Y+���|>:l9��Cn���z�9�-��b���?5�q�_X8J���c��o
�7�?^���� ��K��I�r�V>�q�C�
�k�5u������vC�B/b?�I�-cFݜ�֧�?f��ķ:.��y�汒sn��eR>���b�dd������YZvO�Յ�� f�1*�؇�e@�����Q�tS��("���>I�5d�[G�BIIO�j��T-��3%��Z�orW��q�r|�2�@Y���FQTQ�e��G�Xk�{�8(�+x���Z��jb��c�H5�o����e�њ�Y�=�$���"쨡�����,��@L�'2���(�$+3?���c��\��_�sn����ژ��B�(��*����y��͢@ݙ|Y�+�ۍ�C�PF�F��5,�N
�5�������bY�VxҢ�Tޤ�Z�j�]���J�vv�+�B^Y1;����)amլ�C���Y¯�����~u'+[[����������B)��_����V���#?�S22~�^���sY)�֬�f���
YSn�d{yh(^�1��'\F��ϗ
6���vq� �k��"T�Do��ih[MqLSDv5�>�P���8���r�JG�%6�f�ş@�0A�$�����n��+��mAK��!��J��?�;�
���ő�RSYy�p48O�����u��p�>�k�4��Z��35u6u������i��ḁ֞}�R�ۤ�I���O�/���Zd6#Y=Ȉ���8%�4(�Zv`᜚���5���G�g��w�;��t�\dE셦�0��f���>����<�TV$�:=6G����� ��`�g��ߢ�����'�J�o�5�o�Q�����G�W<����L}�6��4g1�
�[�@��KR��iEo�����M��:�6z`��:�%��\��-M��k��1�m���x���|�bu�z�LZ�y��hnm�E�B���S�������� ,� ����y#��]��>[RR�a�	r[���>~��os��8p�9PX����z��W;����K�Q.�L �:;��V��~�[��@&>=��_���nD/
}���^�i�G)��K~�K{|�!i��yT�j=#��
7�G�G�U�e��S��?�N�> �p������?~Zhh���M�fpRZ0��\\��3'����h?(��)%+�n,0itAEn� ��
{��mȃ�dY�5J�����Ƚ{m	���K~�܁>�U�y��J�Mb�y�Vp��Kռ2��l�i�i%���$,�9�F���L�O��H�J��2�<���=,#�hQ���u�3~8#h�������Lړ��ee@v'�6�H6����Ҽ� ���&�⛛��7q���M�ʳ܍�j�fY��V�h^9k	@@�W�x���)D�!f@�?�@ y6�J�~{t����{9��;�a�;�}��?t@�HjM^*�%)q$�l�m�_y��#��X2݌*���΃܋ћ*�(o��=;���3��n@��Ƌ���G&��ask�i�n�w�����Vi9���/�Δ���E{�,�ǧ}�=�!�;gg�Opz�6�uV:��mvɅ`"Ћb�e>^Xpގjv��.=�1��!�|<=��YE��9k�J��E�;7hy�2�����,O�ru�+��V4�ܚ�ݝ�?78-�,w:�\	�ѝ�f�O���.25��r��݉ VDn�ȇd[��_6#��}�	�w�bo���dcA�Z]9:9�OVİ���˃!,t(�絡&�v�_Ё�tr"x��- ���> ���W4
~a����hk1�1&����q�N��W��A���,����Y�;R�/�m\��oѷ��5448�>@ѫ�#�u�(�̍B���ל�R�$E���ΉWQY����H�a7ĉ�s�X׹�r'g�M��響��(TT�U{���ee����㌢(�^�~^-����0�$(2�I��D���pLI�&�
�Aqn�6�m�Y�=��6]��HO�奮�����7X"m�H��f���R� �� B
�}!؄�N������ �%���ll�PYL��_�޵�,ȇ�Ʉ<�-'��>�_���������G���@iCE?l����DE�+)�P�AM����bZm�w�؂�N����{�މ+���+�i*�]�ͷx4_.!1�����^�>ŗӳ�aY����.j��"t�{���
1A�P�NVތ�B/�$�h��G�e-�7�/�0����ސIw ��O�M=�n��-�je���	/�I���!�	��EE���L��b�0na֚��8��6<���.#픡��@:(G1E�|���t�'�U`����/LcP���'_.9��_�SC(�cY#-
L<�Wp�R���1��X!��#Yz��Q�	���K�S���x����a��r��V'l�K����Ó���K���퀊#��)�x��e����I�����ᐼF/d����@zh�t%z�m4��g	�M�޾j���
0��i���`d��`��lF�e�(�=܏����4[+T~��vH���%������ة��amm]9������i[�Ċ3�%���^��y}�z��Yqa$mʥ���o
�ֻz_%�&��QL����W�\U�6 �<�"d~�wI�'��E�K������4���|H��6���趁S:���37%--Alg�7�uY�㙘�;J���D8����-Tb�Ti�ka`|vn~�Tͬ�=�do��T���̯��s��*�i��0�o�ש��'��fQ �(3�)�Vo8.����IG�pO0]���0ꜞ��i6��PTV^�'^��S�?7�jD��6!�r̖T�ʰ�2p,7U������h:��},�/�wB�B�����4?�T�!ݤ�,U���d�Z �"�L��,��f�0.O�}�-�������UM���P���ÔG��W,�٪��F�Apoa�<��˦�&S �f��0��ΰq���ZK՟\�j;���O�����9�fB��L�$U��wY�y�O�ĸje ��r#���XzJ�����W;�T�=>[��x�Ѥ�{��>[�~mcV�|KD�YZ�].G����\|�:�er;;eJ��t/�w��UB���M��>�����(�G@eRP�!� ��6
 ޽''n���N0|��ml��.�kr��[��٢�qTZ߮*Q����	2c՟RSS�����u�x)#+[(���LE�%��>Y��\	����jE����^,�Ŀ��())�w�%�Ť���F�d��qQ�P�K�/a,:�u�������s^��iԼ�---56�!_�^��e�����6g��G��
I��!q�T�u .`dww�PI��{��ss_L����ڰ�n�"����,K�= 3bb�|Q��琞в���oG�s�Ա��ft���+��� /�h|S.���;433��w��T���tM��=ّb�ټ�M��8r�~���Ac���t���� Ea��GE>v���쾱D�짢E�����oI����g��gEG�;i_e���&�׵gG��,� �
�ȍ���<f���/>�o�@�r��Zi�iJxs���.��Ϗ��� }u}������Y��(�ߵ��w�MT��O}s�-3�Eb��]��k w�}V�o\T�4�Ծ��E�*�]��〟���H�z�9>���x� zz���b�dc_;���������ۍ��O����1���]O�>Ъ���R�1 �5�������_�"FK�R��>��[�ڑ�C�b`�_���ܺ��`~��Y��.U귾�X�l���k����L�i���*~� �^�~������	���K��+Ð�(�%G}��؏r���[>OC]!�UArү�- �Z��1����q�1��.5�|u�s���Ҧ�i��٧q�n	I�C������$D����|���W'z&�p��݁.�����k��@4�[�cb^e�Xxy5���!�6�/'���]�7���;:G�x)�榜_����,ll�{�k@h�@��!@`���%��D
��ڧ"�'���)�@�����=N~~~�ܯ��6j<,@}�(P�V@\ǿ�1��O,q,޳#��9�l��P�p�bz��P�������b���wn���R�>�v?3���b�K#~d떘Z�|V ��죟�N�c1"�:r��3-����w����47G!m�Nh4�wH��#��RX3o�X6^�-��M/+����9:��	E�V+�T�W,���֔��ˁ�<'��~����ȋ�#M-����?n�ss]��ɠ�����ST�3Z�~ɋ�r�"��S3S��7�m�̡53��� ��Y�!7���2G�B���Jy1�1wQ��g�%N � �5z�Ϸ��@TU�ޤdҾ��@�ZuɁ���6btc����-��ї��`�M �L�S�#�>t�s���R�!G>p���L��C$TH3��Қ��ᮔ�o�2��4^]vK�PG0P�B����ӯ�)�:^���W��M�8�V�	G]��K�S��Wa���co����7�bK�xR�j�O�C'B*��-x�ب��t�L���]����+䋝 ՝(�	n�12kn�/� �5�$�DYrq5D�<���P=Ҩ�Lڹ����ȸHN>d}*��jsns��h+�����c��Ӗz��d8��3�=_Q����vm�<������U�/�{Z0��У�9���N�? b(@������O�r$�Uj�;a;�X��}��#��֭4.�Av��d/���|D�  
 Tz�q���I�s��('��@�O5�~ӹ���Im�^^�-��/�����'ϕM�������Z�`��A�;C߿@1��~Nr� mޏ���53�U>I�����n#B�ee8_�����쩔���t�������9��o*E��xQ�Գ��gq}�F��{��ߜ6�}pu�Y������3EFt8OMCC���H�B��FUR�ӣ�&��7x�0��?���Υu�X?�I�.�W@YO��O���^vϾ�1�?��4�I�n��щm��5���×�+.��ycO"�<����Bi�~})_\�S}1�6й������?�;�>ׅ
�	Cc�?��p@�w�}�)��3��rmy���:��95�8̅=C++���`��A��d%�Hcn��#�L��4Pu�Z��Q�塞����4}���Q�03o�V��44���rN��.5� /��	�-��o��I���:ѡ���@J���^<]��SW%-d����3U��\���6�����h�A�vM���*'��Fl��ڐu/����gs�v�9�RΫmԃ6W���k��rfY�^�p֛���J=���t*x�}�}G���%xN�=2��N�{O��T�"��)��f��1jF7�P6+4��F٥���d۫A>��x�̥��u}�as��s�Z�m�QQr��{�}�o�f
ϵ�?T� [�o`�Ng�*9mjO�
k�%�s^���2�ҵbl����B��w6��p:we7\ ���|����4f��R�W�8� (���yv� �Ε�L�(&s�i���6u�pg�7������PeP>;���Pq*��\D9�+c�4{
�vj��T�� u��&FYbF!N`�/r�$��CQ�'�͍�#YG���^�J�H.�X�eƘ�X���M��Oa�6�*~�B�z�؊*�0!���:[T.�(�[n�@γ<{��ǿ�ݙΏD���y� ���$[����Z�	o{̉��M=L�bC���H ��_���\5�ٿ�QVa���&X�-��r���?F���%l�4�%B�b�� k�k�g�q�lG�{&�B������߉_0p��~f�n�Q9�վ����M6H�	�M����_U��[��[ɼ[��)#F��P���O+�]�ب�_�Sk�ę�p7X�Ŋ8���!��4��,�M�qtؠx�Hy�X!���Sd�E̢|�J���M����v`��E����#��ץ
j�b��r�x4x�ZC�w���&"3Kv���J>e�t
�G��Y��H��[4wo��9�O׷r�I=���"4d8��ki��zG��T�z_O���[<��%hBɌ�Z��sg��|���i�Ō⪛I�m3���c,x2��>ǎ
�W ξ�����]l�S{�'[b�k�����P�0	��j������A,��Q�l����R��y-o���ט1�4D ���-iᤤ{
 �з@�s�ϞBa�kذZ��9Ŀ��/ď6�I��!ǕF�#>9ȳY�G�S0PU�%%�l������4�^��a���+>��wN��ȫ�_�*���@ӻ[���d�׌�z�O��[c���:ӈ4���:���z�ކX�-�L�9$c�g݃A��tq���cKtіئ�����G�b���.���u�*a:����(��y��ݻ}i�`/��^��o�3�n{9�rժ��li�ܑӑ�m����[��p2��"t}���=���g>��h��+�Y���?����^�������)c?�B����q����|��r�i�N󍐹���zǵ�����5Nu�����a�p��{IHV䂫��@�5��b?��*񾇓���������[[3��r�l7�D��I"-	[> 5:
�3ɘ�����OX�!�~R< �jP�.P������d9���C%���`���do��N������K
��f}��A�=�^аd� 2P�;)��Q���)|Q2i�th0Eu��G���0��1�ĶA[o��#�����Ї]��q���̡�~�( �f�`���_J�g]%�a������д�"���a����6�e6��_R��f�.ǀ&�sw	3��u�çݿ��U�v�j�+�,2�5�������0���	��?�A
�w�3���G�S����x�
�Kѩ�҆��3��w}k*w��� ��P�/25Vk�{��z`���|��Feۿ��BE����-����Z���z���0t�Ej��<�-�СL�>��ǴxD�j-��A������"	MN��F
�奊�#}|�-�-ʰ� ��9ԇs{j޸�B���o0�eg�<���]5|r�.9DEQ��\��������%�v��j���BաS,cK�Z`�n�("�N�{�{�ٕ����8����-;ɥ�D!x1(
[<Y�M���_�y堬���=$�]���[b���*�`17��p��)>�"'Vgܥ�]�vM�g?��,��K �[e�l��+_��������D �FмPl�T�0��-5�af���4� �w�_��J��|�ՀZ�\�aȵ�u
փ�j���Ra"�Ԙ�Y��"I���\{�Z8��Ɲ�mԡ)زq�*k���z,%8��^�	��j*�e���׈7��|mX
�8�������\$�<�V��u����a�B�G��x����Q0g�$����y��S�[�}'��F�n���o!=�GL�=g��B�!6��4��O���~�rū%��������ps~p�F�do�`�dC�!��|;ǈ�0s�I����?y^��BI�w*੄�պ�o��p���#���d�v%1ZjR�9Γ�Ѣ.�A#o��:�/�ڍm0�o�p���
�I��U_�rtn��l�6X�nc����/����`��O����)�C��8�%�%۱W�cr�����!��.�+S����J;*�&���� �8sU��;�Oڿ�ڵ4�����D��)��u��b�A����#$k��㕳M�a�:%���?Fj�}Y��kSm1R�cU9���t��������3I@q��/6�_h,s|���4h���������Ը�S���(O��L�������;.-ڻ�L��4�C/q{~ѩڔ��h���\�c`�Xa�)��7}���*Q#4`)������0���ݬˌ��j���q:���J�C�y�ӷoc"c��[i�/w	��y�9nz3�B��5�{9�kt�8_�ů2Ba5cnG�)Y��>�)OX)V?��q����૿�����ߔs[U��[��%S<a���~c<L���.��c�S�?�I�?���)�1˪���.�¼O]��p�O�Gǋr����f9(���P��� ͷ�@��dÍu���Q�!гߒST4��Z(�q{(.9'7wHj*e��;�K������Z&[�pd
�9�Hj�~��,̖�d�`�	�DEl��	O�H_Hz�`Vp,����n�.��ի1�>] x�k�EN�ݕ�G>(�'��K��K�R�Z����M����;iS/ͽ@�͖��X�c͢�lO��L���!N�����/M-=�
�TJJʵԋ�g�Z�e���RYm��#+��%���n}�*5���\]Ւ�XRY�GLƯ������
�3��&�_]]�$�m���*+�B����]؉v֓�y]H���0�������ɧ��Х|u��I�G��d7�/�}ydȵ�W1U�1i���ОЎ�~_&���9��g4Zf�G��E��1�5�X=��9�<Roj��$f�z�?��R:�E�/#�q��H{���2<Ӓ+H�L�\?���?Z`�SC��߁8R?�⚕�Ĩ�b@c_Cˎל��f�%s�<fw��0en�Xt�o�f��EB.<�&Z-{�2<=Z��NW��F�
*�+W>,6��_ƒ�|�1�&~o7�&�7��=��q31���0��%�k�}%1݅b�g�1�a��������q�}@�˫��<�b-Z7d�T��<���k��ߵ`��~:�;o��g��u�b��'��L����b����F��(�^"�N����{zj'Y�VW�����3~�u4����7M�ʼ��c�޿}�ҕG��b�/ɤ���Їo�|a�q��c}�W(��Q���rm�GETM���͠?��s� /������N����F��@+�M��ѫM��5�W=ߑ����F�A��k�Sṅ{U?�r���#�G�?�T�36�f0S�����{�]��~���1���$H�0WL�q��Eк�7�J��~)�'����;�vJ��f>��w*bqV��j\I��eL���TN��X���lܔ�{��O~3ѓ_��-u�G���N�5(5ޜU5��'ܹ���H/əP����x;�	�����݆�@��E��:��)���A�6c��|��l#ήZ3�)w�΅�ˏ��k��QKJ_>�K�/�l5rttLGl�&����3V�,ĥ��c%"}j��՜��K��<)m�F\|]ݫ�y@5����*4"��xK����U�z���gi^q�ǲ���Ⱦ���Z6��+�`,�GK��^M�X)�$-#K|vn���U��L3N�|1Ϙ�"8�~=�Eg�h�鯢�#�2����\FqUI!�7��b�����j��a)��N��f���h>(F�/�g��(4?)���j�П�D��iZ?�~���C|��|��se��޷�K�����L��6s�EOߠ�s���-�_ "������WW\���MU�+�l��豕 ��xX�۹�wv�M#������k��Wf�?.�/�O_�Q�uN��G��|G������1�|&g��r�3�
v[*0��m5��rS|������D2��]oB�y�����#��m�z$�G�F��=�c&�\\��2q��؟qg�����)�efM7±t���Y.�wZ_�(��V�'o@T>k���{5}�c$Śl�AWY[��̶ ��*� r�5y�S��@�4-#�}ܽ�J+ذ��o�G�H�f�+�<��9TU�!�q+�s�*��	X:���g��: ���Y�?N����(���������9t�ͦ#�����y�O��#�$s3���<�t5�RE�&ĽH$��XƁ!A�e�=8֧F-1�Y����&��N
��隽1�;y�})����1���ڱ0�`��BȈ����4�k]b���N|�f��0&�S�vZ]��a��r?��͠�T��'˨h�`�w��Y��f@��h�?�kvR�7��-�S���u��x�j�	#��L����^bX��,!�Jl�̊�[�S=������q^�T�������1��nz�-�������7�ʟ��V����O8�Y�~�q&W	�R�G��̘?ֿX}�b
�H�E=j'��o���F�P��-L�K�V�z�w�.q�8�}�ݞ~����c3!�m@��0���7�{�r�	�V����B��_L���dK������ԎI�J��5�Ȕc�N��0\�-��׳KN��޽�u�G�-,�K%���\�y(~xO�(Ƴb[����-�FL=�#~O*��k&c�(����$#8�c$B�9V�HXNǎ��?�ji\�\����fiY�T���ҷ���)v���$���|J�����i)�)4+M��M�v�B�B|j�	G��ΰ���`�nh�0x�P�n2��=�BP�T�@��t�h�~��p\C�'�1�}���jށ�A�6�s��| z\�bI�[s�Y�B�Gj�s���u��2m��p�N:��.�4	\7��5��q孭Fc����R�s���lmm�r���H�>ٱ����]\\P�qJ3}�SXp$��kd2���]�ȼ�2b����1�������W�����I/� �����W�BNѓ�Qx��?��\%��'��>>�%Y���EHm�i%`�چ�M����@}J��K0�i�Xrma��<��{�5 �S��6�%���lB����9o4�-c��r�;��8?�Ҙ�fd��{U��P�.�N:�*I�?|�!�,!����Y���ϥFUm֘3��I7.eS���%:'��5=����[��/$ ��F��o����{����ħ�6q����Si�=q��,����'��JI� ~��ȴ�ޚ���R������Y��e� �5|rWL{��"t�����Zd��I��<lU�;
8s��Π�,e�N�(2�<�̎e|-M�qUm�/�����{�6P����[C''�)6_�O��J�u���x]�?w��9�<�35�M��||}�����[���ut�<ycI�&o��ԟ���By/��?��|�6?�ݦ���ڡ@�s�k���� N*���>F�U�v�S٦羆۔;��*؝0w���@b^x�s߼r +�ZL^|��xS��f��G�q2:>P`Ͼ�l�U�sE�:�Z�� �E�����8�l���kؘ�a��<e���H�?w�mg�{l/N%/��o�?7�'��~�O�����e�R/��ȺZ2�6��f�ӑ��d�8ǍXTT8�ez RD�S�b��W?镻�o�H�%�U�e���&����ir9\����p&����y�̶w�0�%����/�RF�$�{"-K��cK����Y iR�d_@E	�x g_�>qBϷ�,~���o�'��P��P�5?���P>�6�]�x�s��)�#�ݝ5�l��q�ل�C#�?��o���F�b����B����#��|P��-k�4��ҙ� xe�2�YYX�����8K�0�ք�=�%s�]�>�ۤ���ѩ#�����Y���ټ$$�7r��o�w�%���6|y� �耙����_���Ͷf7�{V��{klevm�2�\�Қ[�c��8����	��L$V;f4��ic����J7w��M�G�p�:�M�W��vj�:hd�?t�]��y��Y���)Xkrښ�f���iSQ�}ۧŬ�Ͳ$� m�߿I��-ƃ�oi��f�[�[`��!���5Ya������}�V����p�;D�T\;C�0�,�ZZ(�.n�A��+r�yy��/~MG�m@��U"ms��T�e����w���|��|���U_��=���NEG�.BW�o3A2��w]��Z�,����ݤ�z��ل�Uc�#��i�		dɜ����s��:Ԍ��HsG؈�-�=�����R�	�Պ�&�w�3H���~s��/��nYt�?Yc{ۏM:���(7;�ӈ�dj	1=�է�|�ޓ{5�_L���b?Z��.��s.v��d�j��d��)�'#��kx�O��Sj�"@���������*s�	��Ŝڎe�)�߷Lqj�19��d��Ѣ{�H��&f��*l�z�V�Hq���	澹�.�p����Ob^�u�{�q��K����6�{�c�O�m�a.j�|����o�+[�K�;���v�����i�����U�,8�[��p�#�o��7x�;�(ߕOٗ�6��	F#˔�H)����z�1�-a�0� Z������ ��#F�^�0���9�"��ʍÜ���8�8;�(:�_�����3/&����FO&�S�* �T�8���/���=�>T��#���Q���lI�1��ܥ7���X��`���.f:���i�Y{K��VK���9�L����z.��ɴS���_U�G��ϓ�+a~�E~��s��;���Y�q�4�V>��v�v��+��QM@M�Z��J��3���K�sXG��o�ۍ��C�f���a���e��YXIA����/�O�Af�#2\=*(��]�����S�9�2����'k$s��W,g�/>��mJ���JrvŘGu��	׆B�++�KwJY�k�9zi���_�u|��D<��O���J���P��K�_ 	$�SX�o����v���* �$����>�a]�,���-�<�.������M��4�@�X�AÉH�����E�;!�׍[5�_d��p^��s�@#��6}d��מ����8�����c�R/�"JӚ��U��Rl�Q���^�&#������<�d���:Q�f�o9�ܳb��+'2R��p���v��XF_8~���}$T��y��qC���SDg��E���N���J�L���}Ο)F��W��?�0�!�Z�5خ�'�sl��������C1��	�D�[1$�JX�Բ��J���FM�l��y�tDK�Z4ꇦ�����c��1y�(�b\����u���6�_�;�����-v�O�$F���|]I�*9�FgT���x���!Y\��S��tԢ�f�g үI�FK�?��K���E��2���8�8�+��B��>:0�ۏ�U�a8�����B�>����\z�_�;�Ð��@�m`�]IՁ��i���z�f�qK	}�DPP^�%~��Ω׵�6x*��2�Ǖ�/*q��/���]�`�V�9�B������T�t"�"z�Q4��'����O�;�
����!��ݤE9x�����8���E�,ϳᇒű�7���S�Y���1�8x*��4R(J�����5L����j�{�̉�K
�g�œ��G�}��L�I�m�q��O8�.��B�9�+�y��<�T��=;H{;�ϼ�	��8R��L��ל?�dq K=烘�t��t��g�Uz*�)S�,�[�B�
*R�ԑ����k�^�"���7�[僲<{I=�r�3���/���a47�,�}���{?�;�7�~fx�B ]?+�nS���Z�����,�++�@�f'�G%JB��;��ĳ<�@iU*�Jx\��Ǧ��,f`>jx��[m���-�b7U��=i��v^$t��2�#>7=� ��T��hD��yyt�u��_F����gC"|�b�;�+{Bi��W2��c@�d�����<��_"����Z�Uҝ_�ɸ����&�t�k���٥�����,k9k����k_��sI���>��F2�������M���O�Hŧ���|�Нz�v���&r<���w��Lm���2����2AߩO݆��Ⱥ�U}eĳ���*=�{J�H��^K�F�!6��RN�����Ǌ(4vf�_l�����6B�����n�����m�c��}��yY��g.��.���Op��{	2$��˿��E��@��T5_Iȸl+�@_FI@��4�� 2��%�fu�vq�d��w/��^4���{]�?E�;-��px��<�X3��}X����ZB��o��⏺Og���/���w��;,
�O ���͌��|:�|*;�)s��[r��ҫ���c9p	�E�"@T���`	���4qbu�(lM4zLX|C�j�̋ί��?�p�iƮ�/X���s�Ÿ7$9�|�����e�f�~��߫Mͤ@67�EW3�s��a6�k�tN9�I�n��Cn�/�B���<�{���r�]��@ͥS�N)Z��S"xl�w�RG<���V�`�R�
=Rpd�X� D��F�y&;��������:+�;|S�,�\B������ڞc+Qk+^=VE�+Z���(�������q6�����	���;���P�o%��r������Y�������ƿuh-����:�X�9C���d^5 ��=dϪ ��,Z���U�3d���qj�Mp��8 ����J^&3�VЄp�6CH�hӿ5���k�/�ٟLOc :�0����IW۔�Y��NbC��aCk�ɿ���O��ۑ�����3��[��iX凓��6���~c$�A��J��4�	��u�O\p8U*+��8�v����#��X9U\+����������!h!m�-&���H�/�!��ˍ]r��E˹�����'��@([���W����.�ّO���{����f���r5���|tQ��Ȯ�j
Ѻ�������q;�&����� ܤ��������q��L!�K{3m��%���\�ߔ�����F�w	{P�jjEu�������0�i.T��履���4oe��u��Ev@X�KCi��P�$@V��2#vz%N��{��`�3�Q����^8E츽i�]2�ʿ
C�-8>I
��8W���2kkj>�r�*�F8�������{&N_�k_ׂg_���p ��[�FK�c���٤�j��Ty�* i	6�q����s�!�*S^3@eF�7��ا�G��/�@	i׉Cq޾^R���>�e�$�;2�m��Z3�Q�(r��;�ʔ�B�������'Z�/� pM��8�ތ�Y��y3�F���b�6s��׎A*��ja�_���чt<���s�&i�u,}��z�bͤ�*��C�i�C7в��DFszA��eg���?!h���	Y&'�	��N���Pe�c_h�jan;�aC*X��~X��͋mӎ�,>~鳰���I*�2#����#��S]�W�\��#ҭ*E�����B�I�+v�����Ay6��(��Y��]�MAW��
��P
a��;���D��K rE|<׊�hߏ���$*������f�2.�	9��dd_����:�2��iWF���h�1%k��خ��ɶs\Ɉp���(�voT@���0���3��)J�.W�)� ��WdJ�2BZ8g�	� n�=!ͣ�S���?�}&,
�dM{�Ы ���9s���B��?�1��]���wڮ����"�ƢSE|��MNP#MoLFدw���r���vo+0�*,��խ���i vǲ�W�Q}��s��6o a��o��fK:1��D�i,��G�����сS��T�1n_>�iN#k�/rTo1�:�Te�E�S7�K�d%����O���3��JAO�CH�	X������O�. ��H��(��%XE0=c�bE��2�E#��Z;(ϣ�3��%=v^���'s�(5v$�Z(��?v=5h��t�0�����Q�F��a*��I��ۨ4�2ش�
�n,l��b���׽m�5�]	i�mG���*Ȭ���1���Z�*s�)'/(��8��˧s���p�V[����������i����"�_i�	x����o��NE\�o7V�f�{��S	���H=�������®�����
�~*9�Z}���L�*�3�[��_N,�<Ǻ7��?�C�k��vX2�y�Ǜ-�0��OՀ��ǳ.�^����Hu���5j���<��$�	�%����	�	 ��]�w,�����{�{7������3E1�ݟ����^�Ti�.7��F�vm����c��}b��`�^�����eے�)�,cQ8�yD�F�I����3�m�4�)��Zh�n�OP�5W˫�Ge����EԮI��O�C"}�!�5� vA�baD�i��g��vԜNp�K��|�8eΨ�ǆM_(,��&�Eq��mg[�:�Z[�M�ʧ�� �6|��˵gR�
J-�h�6��/(ޑ��L�|=�Br�����p��n�6��^�c3����4�/s�3�@3�Jq�4�hn�nZs�#2�0z�t�9��>��O���r�!��%̜u'�L��	�%?E�?fi������՞cPGOtg��K!�/�
�E뷋��E��~6C�+���L�T��<S��]�aU�����C�+��I�n�Wg&m�j}2Q�7��|��y�A�h`/�F�6-�1�/�|j�IѪ�*�7��<�H`Ń�o�g.r魭@��?l��1U^�k���ҽ7�9��9"iK��5�fv�f��W����#�&��K�`E	|�JQ��m��5_�g!�#��9=Y]r$�+ٛ��-r���a�~�h"ls-&=;1S*�Y.uuߕ�OU��:�m����u�|�y�o�T�f�xu?�=>j����咦j�Dh��Ɗ�g��U��3�`\&cy!��m�Hه��l�u8)+M9�#�؉Z���6�����NM�Y�6&���%MIM��*\�GK���S�\��5 �c�]��-���d:��{���S=K������"[��&��R��W5�Ki{Y��kYz�l������-���S	��B�ɭ.�d�R�I�j�����R�����2x�'Z@�߭|��"��$�F4B;�Xf�ox�*��A��&��/gW\���8v��ܨ�|��oН�վ5�0~���"!���SoJ����+�s���1|E�C�**k"׃w�������:�M��b�C9X�:��]6]i���,���ۢ�����������������J��'�S�&���ͬ)5�H��Y�����]zkE�^�3#Vմ�f�8�k��Z2�H!@T��2�W ��������IG�I�는^j|ܙΔdL��O�1a�
�ߙ�XV=�O�)e�w�V� �<��+>�Twʱ?uuD�uu���I6Ǆc7Y��C?��r�a6�}���w�FQ6ʧ:�4���<ܱoé$�!hcl4[�(��l4�D�+��	�=�$Wwf�$��3�K}���ۚ��`�*��.`�������茭�j�1�
� гU��U[�i&VQ�0P��2bI6{ֺ�ȍ��ʕ}����HJ���ݗB��y��v��Q
�d`]}u|�L�́W�Sߣ~u��O����KC��Q��?�A��&��� �� �%���i���r����7(�����]nv���ی���F�c|g�} �g*����C��:�PZv��5�z�W��9���Sa'�sa�j�Ɔ�bx���/@�]���:?ܵ	_p�\���%@]x:H��"�s,�m^�+|ͺ �u�W�X���f3٧��	K�:Q�尖ŋ1����/1�W��7Ժ�t�cD���V��:�?N�WN�=����9��Ar�/�v�}�v�϶�n�6�F�c��M�_� �)�]U����,@���5�ܸ�Mbm����
�ے8�#x�����ǭG�9w�?����@���:,$���%I�a$����<T�3�����E���+M�]��K��}����w���]bWO��X#�Q��N�2��z��xc�_����j���M��a����p�~�Ղ][�U�V%D��i����gWoy;������dF���2}y��f���A������U��7���f�E�XeW�/+/Q�w:ڶ�\��n���v�V(ِ\i�j�o�d��8s|O���Ps��L���!���0L�D��ZU� J��w�����f����5�Ѵ��V~Yc;�|=�Q�8�mY�/��i��G���N@99Y�g�Ӂ��^����@ݟ�J'�a��βzk�Q��x&�>�es�A�	�x+�7�.";A��g��(�k;'�F��<�~��'�{�}(�Q��)N��Q����qh���h6
�[z^v��:�]U��c��l���ɀ����E�ͥWY�8��I���)G���W��Z���
�����/���&(�o����S�n��Z��;��������ĩ:�'���%WU�8�Yu�J.����I���h������a)���K�k�RA��R��u�2���)yby���).�ߵ}\�T���'���y��ڵv�����	'oW���zZY���\���="��l�����<��fw��@u�WR�::��������+Q 6ҝdFM�2O�|"��7�F��<�ד��m<J}U�sp��e��^q��<�|"rc?�O����mS��u���H�<���;=^}a^bb���(�����5����K(L���L������!����?���"����^�@0�=��í3�L��!;�׋6�w�����������4u�� 0�?�H��B���/. �"������,��?�~��xi'�����9,A��	���]��i��4s�K
�c���n(Ԝ5�1�|3���%9�;�n�E�jk���Hi���NNS��Io��]J$��%��x�6��Es>��$6�3�=��=�:J��5�u)�1�B1�UL��5u�Ώ<|l��h�q҆�#"���M� ��T3�L�^%��k�{�D���J,�1�oG�R*b�F~��l6��낥�ח�5M>0���m]Q^��F�P���|��LZ;�H/������|�H\����ڡխ�Z8m���
lZ*�˜�^!����5}���MA����q�OZ�o����g2Ҧ��h��1
�Q�����S̥.��gq.����'��
o��s������WJ�DY��ҷ����~S��s�k
�OY��&�jC�V��u�8�=�/��nf���Q�HU�]Ĺ��ɒ��b�bH�eǓȿiԭ�mJoc ��m���ΰ'�y_�+�շ�k���4@��8�_�<��^���t�tY� æ�#C5�.���_h���E[���E[vD_����@ciSoe8�����C[K9B1�zN�-+�u5_��ݞ=�/Xd�|cy�$�z5�w���}�?�l(�޽��ǽ�R>5�nbj�e��U)�|x�S�?E}��Ǒ�]n���/ۧ������M!b�tዱ8K�w����ܵ&�q�=����)0Bؗ��e����*��TQݐ�d�v�y���[E֟��A@��/I�u8D���nq-Gr6�g��gx1Q$n�*Rcz�_�.-.D)$* @1��� w+cT<�U{�L��CD��;��6*��>V�����J����?r�̼b�L"o�۵̉V���.aK�����S�c���4�j����;u9�0�/ny���Ι��d+%���Cp]�SE�s�U$}� w��ҕ�-�A�<2)�&�~���hk��W�B$���@�5�2fсT�~�y?�7��
X��p���W��E�	a��+��P���x���.́����@�Rl 4~���G�4j�?<f�<䨹L#�tʚnW	9��F��c�XƑHޞ8��)G"	�q37�<��D�&M�xS���0��"66-,��p|�~�4J����X����\y�ŉ�c�2kEb�	wC,��G3�-rT:u'�w܏�����6yf�X*�ӏV�/|�-U���Y�u(�V϶y�SK����K���A�Hi�˟n,D�/��I�G���������*�6�nj������P蔏�C�
Ћ�jq/u��ΏԬ����?������9��W�/�9$8���M<��Lm�.���rֈ46��.���$`+��n�@�X)�vs1T�IelB�6�?ݿY��k}���]E�q��λ�p�2��v��J�	D~.���`�7��?K�F�"@_S��s4?���)��邡���;�2�\`Sy��H�rT�	$�\��f�lf�ir%8/�ȡ����c"(/���������v�&�Àh w/c;,�mRx��������Um�������bcX1J�%�H�F��;�i��i?�A��ϳI@���nr�(�g*y�،��5�݀�(�j��G�_�d#,����#�Y9#L�,��q;�ɾ��Dt�s�|p˃%>���+�p�.&. �BPp's��tF	�ťeeXMN�﫺�����M=��,Q����f5�#����Z�
b��@)��Y؋����3�\>�~���K 1{plp3�i'f�����Y`�ټ��������ͥ����̯�-�/U�J�q�����ֲ�����<��^f�����i'"�a�s��6�I��k8*����%%fy2J���j�b"�|V��hRL�����R3�_y�'@�(P��T*ց	�F�>�Vz�[��"�t�Yr�T+$�������$
3�_�.�,�O?kqǇ4q�4F�1����D��g�����^9����
�?�L٢�~��V�^s��ǡb��^���8K ��}�(Ͻ���i4��|ӽ����,o�JH0l�)������K/��A=J�ܗBCJ1{�:qx�{o��n�𼉽̨�	wh�#��!i�K+����`1 ���MpM?U�be1�N��I���Sȼ\ ٌϓ"`�&゗�ьƀ%�����F�;��X&% 4q�jF�.��?�xK�-�*����B�0k#)�z5 �W�e��<^ �6�k�D/�#����1El ��'���L5��@Wc�nW./v}�4r���8	�@sР��%B7:a��X�^嘽��~Ѥ
_;�'���v�oL\��)�����x�R1ǳ�0{��_��X2<�R`FD~�5b�*�V�0I���T��u��$�0�<�WsM�5	u�UζG��s�0�0k�@3����EL��ξx;��w��{�r�<�T�:9m� k׎w���ek�ҳ����6o�T�J����FI'�nᖛ2d���W;lzrz���vo���%3�!uV����eIr�}�^8Kh�;d�2<�U��1ѻ�T �4���vÓKEJ+>e+��//%�����w�$�}&���#�"����o�" *ʳE����m��]$y�V��5�g�r��4����zSR�%3����Zݶ�z�mb�[dJ�.��@6���72���`V
��6�Mᆂ䲙j���]��%щ�2��*̣--Q���J�Z�c�U.�_�[��@�|&��>�]4�a�zH�DȻ�|��|:��mq��џ`V���B��bb�9���M@PX̬�@;��&���=Ey{کL+{�#п#z0��J���E�[3�0˧=�-T��zl�&����X���m�	(�ݺ�}��8��.I6�!̼��V�k�ߥ.�cdu���?D��V߶;�-��K|��k�;J�![gU��T�
�x���Z<};�)2��:Fy�pD��"�A�v`�)�ݥ��a9b��8r�w�U����-��v��c�gQ=k�x���AxɎ�"��VN!1���O��vu*)�Z�>��m���-�P�������[���� �[B[�i@������<��Ȓ����J �h-��j��~�l*��&�P�ڈ����Ã�`q���o	�,���E�ۛx�0������a+�0�.��Kll�6���Ba8}S�VV��7��%J��M8����N�CNHI��t 3�l.�rf�+yr��@;�9���o�"���J��d�紫*隼?��Ҟ�#���QM��sk���� ��,�0 0�w��^�P��BB�P0�%�d�Qi �����(�f1��L�в��wH�7��U�`4�x3.?�c-��S#�5�?�yZԈ��VɆ�������\D �����g����!ƗD���ɧ
!���Y�:l:�Q�1�m6;R|N�E�RI��õ���}�v�yY���	��3|�c�B� ����*��aw��kY仿{%�|֭�� N�������B�aN80�b�Q��rEǛ����f�fӎl����wM����Z��<�3��$�%�;e^gu�$�j/�sV/`�cc�u�(�1��r�6f-��0ק�
6���@��VH���V/�[|{:�<�V�o�B|��'� ��\��5Y����q)���|��g�ۮ�p�$x���ͷ��\Lo/��|����Oܥa�"z�	�����w�P��j0(�m�;o�Zh��=~��ٿS"�.ݪ���i�<�*Ju��Uׅ���"S,w�C��nO+�����G���@ �1���y���K+yg-v���Q`��a��_����i��(��vp�_ݹ�Z�o8v���2<P�:�&���A�4jW�jN�YD��:�/�}wS��F5|�+�c�_�bg����~����������� Z8�ȄE�� ��]��z5Y��1֓芌B�k㞋K�N���"ɪeOHB���B�i��ȍ$��������	����f�Al�OWMB�L��̢�V�w��Ja�"�d�n�q�jȆ-\s�Ss��e�E;�
�����Q�r�g��\�qy�w�d��_W����?�Ӌ!4��1`����*+Id�2��~���bA[Q��9�/�lsV��ahT_1hQu�7P����!��=C��:�j�?�&ۗ�X?�G�o/�E�a��?�è���K���fN�V��y�/��v�Ja�we�h|�S�v�\��DU۟ƍU�����o���m�����CN�5��-_�8����s!(�Pу,���/j�:y�FlǫkX�K<a�Л�w�&gh�k�j�-�l!>z�նӗ>w���K�#�C'?s�P����$�#��
��(��{lnn�є��׉	�����dEk3	F[�szh�&[�w�H*$j1%\�ҬOq3\�'y�s�3�\�>_I��^''�'|���*��l1�QU��!'�)�	�͍�u����{���y^ʷ|�Cg>�|m.Z��0��|c!Ԍ�Ί� �����fp��-�/��o ���J�CQ0i�K8� ʏ��"4��(�8������|lI������]�� �쓅;��ys�w���﹠��
G�y��09~k��_������V�!'ᨼZ7���L��4�����	��M��χ Jqz����񴜩4��SR		F9\8�o�,S���8т���=�9K��m%�mH!o�S����n�+3�%�mEqP�X�#���F�U3���8��w��>�z,����̢���^}�SK"Q0$�FF�LB%D1�	&�A�����������K�Lt�<,���柑�j����Z�?B�j�t��y���uR���j �RwW+�7J4�y37j�J�nbvI�Ϯf�P-���~��*�B���[�둗^YC�\�����{�&`=A�� ���(�[�so��瞭�G{�i���nL*�;���l_������T\��9��jN��R�YM՜e�߻�y��~��*M5��" �B���<>���-�2Ƚs��h=����A2s��w���`}���^�o^�X�;��t��jK)9��s��w
Q�f�����1R~2F���d�k&���oG�(ŵƞmu 0žw�Rj�s��9�+E���@��~���B�9�y|mʷIT�$����[�G�P�W������j�C\�m.��0��N���w����L\R��]�oM˴�N1��j(
�Y�xvG�_,��K��`��&F�W���>u�EVRJl���:.��F��K�����myk� �%�})-7�:ڕ�Bz	I�p�8"��W��WZK�0�4_BT�ώ.�z@��}=w=y�����)�~�tƁ�l#�n#Gh#�dXw���j��-�	���n��}ގ���Eo��%T0�`n� h_�)	mކ�g�͵�W���Q���S���3l�7%4		�{]^��Jc�M���&A	+cV9��f�Z Ac��GdR�o�X~��-�(YF�z��Ҷ_w��s� �;�KZ��h��\$V�Õ�9!���D��k�ϼ(p@
4D�vo�PD`!�l�8�:n�Q�`i�obi��y@3���^ԡ��'3d��r�����ʥ�x��ǣ�6����8��D��fX�-�m�������
R#?�G�G�*yv>�Ѻ�f=	.�kv.�sҝ���ÿ��>1��v)��!�!v�5�W�j��ЌeZ]M���c�]ea��ߩ��^�����_G.�"��I�r0�z�O&����IVm.��rV�q��v��Sz���vW���F��d��i�Wp\D�\|,B�so8�Z�y�D1(A3�fp0�$�F�\]3���xH	�*��� r^f��X���~,iq����Y�E���i�� �y7�����;��j�"��A����l�%�9l�5*Bpnf��v��!pI�ˣ��X6������E�;���z������2�<�h��C	#4���vr�����v4@�B���e�3�P/uF���A��;���M�_�)�������_��e�&�l�*2�����ɜ��>!92uP�����w�>eg�}L��5����k̺UcS�qYg�B����uG��[��tԦ����=�0�����=��T��y�5��HhS]��'�Ʒ0��k�|�j7��OÆ{-���x�.$h��zvOBr��h�Jt���+i:6�ARxm�B�X��iT:��u�fkE�)eu5�z�M_�Ǒ�t�o��}E��ZH\i�vC�A'��L?�B��]3��,(a���q�i�GA݊K�AG���y��$!~�2�bR�^�)��4���2�r����҅b�+�o�y��y��ti~���2F�\� \�ǯ�{�A�P���������u����6������M �n����[Ȑ�~�f�'M3���k̛�)-	�e=o"��k-��d��E��o�љ�������u�G(T��D��(#.ف�=cޏ��Kc԰��b͠����eK�ݗ�wwQ���s��U�w�y�b�'ح�G,2|6O��(���q�/*����^��ta2-���߄H������릚��Բ0�/l�������������m(�@�~�T~�Dp�,Y]�^�z�ŴC����K"S���K\��r��Y��h��=��0q�Q5���:�̍��|_��d�� [L�z�f�ThV�o�m�^@ou=bi�P8m�E�9^�3i��꧙��2�����+��2�}��n������K6���q:"���ƽ���)���u^�R_�y�5y�?�R��f4�����c<{4zm�t��i6����51�v\�.�Z,*�X�X�Q�Ѩߴ����B���;^`MO��2b�>�1�&��k\.$�7���0~�t���U<Ǩ}�L�����uw�<`9��uL<s���fykp/+R'���
�G+���F�H҆�#li�-�x�M��ā�7D�%�
�s����"@�HI-�Ύy���
6���w�k�Ҋ�k�n�;#r^����}L�uW4r���IN�ԣ��H�<���~����ro!_2TSy��%���"l�S�����/��8a!�>9�S��Vވ�R0��X�A�������!_������k���?�`7=��dk/�p�>]"A}�s�I�o���NNƯ���������>C4�������K��.���˚5�1�1�8<Q�W.��� ���T��c�������@�lޓ܈�tF?a�]����9�g��2��~I����m�Y{���c��i=mj`O����v����e'0/�y>��^/m���[�&|^ZZR,�a;��:��=���B�#���Ë��3�.�:7�W!���鳃�ɚj�z��ˬ�Pl���^�

�vc���:�V�W�C����Q�u&%�" ��2�c�����Jb����J1󇁔
A�8�[�һ����]�9�����&B��;�O%)EI_S9����P��&7=Ġ���`SRX3 �a9 P���6�Z�5�l��s��C��அ����^�����~��%��ǆ�KF1�s�e�M�Qc�4�G���/���%��?0�c�W�Q6�#݀�ؘ�FHcr2��8W�<��� �y� ��w�k3���ya�E���-oa��8Lo]�s����^~�Y��� �tS�/H.`l���Gn��m;�1���޺��SG��ް�"�'�@�Q'F�T���C��4�a�H��wq΂���e(����.�=����	W�79�4Z�+*�u7-���:��:��s�j��{�gM����L�8�۫������AA��d8�VdG�Wyˆ�~�n^�X����gO'��D��LD���R�hx�M����p�3�zd�g�e�ʈ*t�\w?�-&v�h�םFo��ʳ��LH9�욁�&l)�z��e�\܅C����$C#qm���8�]G�~&:�^'������j&�>m@���p�<����a�$\!r�+x;�*���K� >V�<�,��3�$���i<���v�����cĤ�<�܀'�opC�ڄS�gYe�ߣME�@�l��M�$ǯ���>FY����P��ꅪ5<��5��y�M�a��Q�"��0�oha�ol�����������`!m-2�}�w�\���.�s���E�FG����(#�_KT�!��,&"7� �k4ǆ�2�>��cU,�����5U����ϑ`EM�9�.#L�
�LV�/�(my�o��w�$	u��*3@�k�#{!���1��W���8���	���m���OR<]��d�{@mmZ�쟢�B2R*��#��	����R�PR��nʮ1���j��~x�����zﬦ�\�da�q�!���5W�}� �4�J��on�t�R��'�\A*����e@�����bM�a ��-���9���v���='}����T����N��*����k�.h�Ky��0~>��I���W�'�oN�U�(�%�N˰���������Liܒ{ε���.<�	i	\ٲx��|��&��1���Rtz����a=��
u�p�x�ʫ4��t`�	��HO�}7���<�|��Nh����|�c��y������ʅCd��jԊ9�챔ʨ���C&�`@�I�I7
Y�|��y��ܖ��p��yz��U�byf:��x���*Z�	���}��lB|rrXn�p�NiJ�~̤�@�[���z�z��ؼ�yc�>�m߹��܈��^��G/�����N�o9WI�6�������ox&�*��7B��Ϸ3�n�$��0��zT�d��c�	���Ώ���q�I;A~NNJj���:R�p#��B���/��?�~�P���~V	�J��z[Z������d� T`������s��m ���b�A|�6���,��Ϻj0�ͮ���m� �mJ<֍"��L�O�3T(�.�Jd~ʍ�o|��/��+k��C�_�E�!4���')Gv}vy�c��Q ��V!Em��OG�9�FDhҙ�Z�>Tw�7Pn��L5����G���]��%*E��ͳ���鐭-�F=VW����@��d�A��S���b�ǒ�ے[��a)�x�@E����H�[�.e�z��D�e�6{9n���x�����m��{ޖ�0F��c.�kLLT,$�5`ť%�,8h++sfv�j枙��Ϻ�gT�l���D�mդJJ"���;E5�PX�˛���S�I�~폵ɤ�"a��@�3�҆
`�At���1���"��)�D��$�D�ϻ��w���eL�31#I(�>)hJ�f�?I�bm� Iv�q�d-3;���P�_G�������P�aQ������-:�kwR$�^�xJ"�n@�'���2��:�
|u���9F9l;�?� p��Z�O�8[=V���v�a �����2d
.�L�(WG[ʲhXK�~v|x�4g�f�9��S��w���B�n�L�b�N��&221{{>`�o�~m�MW�#�ſ�C����
 j�h�g������C}l����ǡ��"o�^@F�ψTOl�`h��7�n����{{�_D}�����7�9�9��Ā�kW#BE���{�I�xB�,P)���?N��&)b��|�e}MC�"��GH���䱵����z���r�v`p0�ׄ�Eu�%�M0�-�W�\Tl,���!*zLƺ��ro���\�}�K#��KZ�������s�2EB���u�R~Ӈ�L���e��nq�_���n��H.�Ԕ��!��L�G���Z�����&�;`��X���tf�JM
�C"���K@��,o�TK�_o @)����SSy YYK8F�g����@d%�y�aɅ�ϐ�=.�?�j�s�[q��s�zik�m�oN�i�zx���>���D��a>R�����:�˵�5զ	3�Εҩ���Λ���r �eJ��s`���2��%q�q�+�hh���*N��-1���+���:!ڳfF���I�|n�R�����Ȱ������D-�75�=<9��.�&=�� %�iRbMf���#���B��I��˻�`ǨW�b�lX#��t�]U���j����r��?h�{�*���b�{-��KBLB211���R�]��2jiw$�y��ڰa;h"������{�g!,Ze'��>���H������������4l�*Z�a1���5F�_'6W�
�Lq���^�]y|w�G�R����Ģ�6��baBL���9dd�����JSb�Hd��!��z�=͓�e��DjJ���W�ۈO����#���� ��og��KU�.ƴ	�3`ڻ�ƈњ��i� q:)�>�wH�D_@Jzt!�1�_벙���ѓI>��z�&{=�Wҧ�7�f��MZ)�4�|T��� �����|�!�1#=�o�!�Т٧.�뗸ԑ0����O�� �`I��B��`!=M`�{�#����Iѳ��4;�a��Q���wLL�|�EzF���؞����'��L����&�h>:�,m*c^�H;l�����	.K; �@IO��e�3��%��3"�`
� fX\\�Yk�Dr��@Mτ����#���S*O�#՞�:�����Ǟ)�/�+F�y��ԡt�	�����{��.��N6{7/�t~�0$�R>o�tf�{EM��EtT�h�SB����[�gj"���C�#3tb��B8_s$���^�Uм���:\�2�Q}j���ʵ_5P��qZҧ����.��f��B4�+�7�(�xֺ4��*�2�<*�m$$�d��^(J�&�BG�l:�'Tc��wiJX�̓��?!D`5�P��N7�
�^�
�	�8*r���u�\���e����������k3�[�R��w��������t�/���4�uwh�fID�X����S�����Mf16pVff�ͬ���w@��Y����Efm���.��n��>�%>Kj\�/�F��q���A���t,�Wܴ/a	__�]��y��tU�t�I�X2�A�Xe"CO�'m�f8ZW�]��%јX�z1�n`Pb�����6�iG{��&T�孊���{hHu{[&b�Ɣ�̾��G���*&��KK#�N&r�	6JOm��2b��aҦ��V�2��X���]{o�c	�Ƨ�4�^�Z_OGPuM����C�r:��+B9��/Wf�iʪ�A`0X"��s��8�((***���]��\\�[ݛ�-GdSs���?��� :7}�� f��n����H�.7�*ȋ��l[*�_9� #1ΪȐ%�lmN}��À��b��g2W���F=���wUӋ���w~��.-ށe˥�Q�h��[�� �J���=����2�� 5I�'R�2��+�����m�wd}�0T)�M|�D��5���"T�̱&��7�qTGt�)L���<�ŷX�K�}G��]^A���=|�k�A�"�U��q����Cg*ܼY����q�^��͡$~iqq1�ЯS��B|��Ḩ��?�3�h<�=�W�e/�"��TГ���fW�:�_��h�{�!��qx�{�*3�I�Ĝ�s�)�����D�}�]:�����W�}�������GM
s������t����q�Π��������<�)̿b�ˮb�L�H/�_���ey�W������������d��(|�H�ǫz�jg�r�����r�A�3�k�K999e55ܫ�ۻ;���=g�u�ט쾷���B���2���8��q��'*إ룩g[���;��Fy�ǝ�X�����).�U���j��{�%����,�jǦ�yåh.���e_��r�s�=}����ˇ����4<�v����� ѩ�@���?;���k�q�}�^ .N�+�����c+��,3S?|s3!v��@�p<�6t+�ITA�k�'��ע��2}��Ɉ�dE��{��o/�&��&�L*͆�]����#Nn|,��5Z�Cp�:�c��Dl;gB���6rQ4QC�he� �T��V�هF3����;��w�-�z��!J���"��WW����[��U�0�>��>n��a��A__�:v`�zާ�w�ʃ-��e�]4��!�R����[�� �1�s[��������n ��7��Ӈ �;��a�(�o�
{&�-�u���
n��q�[���2}�<�?1k�Y�O��Vf�����` ���'��@�Eè�7W�I��F����!���%%L]�ԘH��H��Ro��^�8���nAT"�-N�zW)��e�y�9l�`��Ҵ`�W�^�x����5�~�����r\�(Z���|�3,,Y��c��ĳH^�ň��Qw�e1�������;an�*Q�ãF6^h��˲�j�U��'���ƅb7���@A���"y��^�\���U�o�D(���¥1F\Ǌ�HrG��_�}�H���_����)*�dG��x0@x6�.L���ӹt9�"��4��_�J=�����.���lK
%e��
Se2��Q$TH/��:(*�.u��|�,n�9a��9��|���f��k[;�U?{���� �I����ag?�I����h��DmB	07�<�ЃG��E��c�ӽ�����׎��h��z���~�x��ު��_�_��VQX�T��`���!5�XZ�=���_��[$�w�|zs}���)�<�6��γ�Tp0��������6e�I��O��/&�F)�xT|0����|#v[���ܯl8��V�y~�X�����X�:d�O鮂d��;���ۣ� [+8Jr�k|�ދĻ�6|&���V��UoKD��^��b���t�Yj	��)?I��;8�9�o��B�a&P7`�ܢm����̄ϚH�9�Лa u��rV�ڬ�hs�l^{9`y�b�%�I���� �P�Yg�7�o�`�R���2����v{}�U��;�����c���6�^�/,�}���`��+¡��=u�eT�}C�gj|���92l��*g
���}�Z���q��C�h�����`^�%��|TE�E���t��[�xBW����LI�=������1iss��ay�σ!����9�H�-hM�R�|)]��[gA��Z���fi4�%>/C�l�gO�-�_�̦f1���ߴ ��j��Fx�#x�7X��8����iב_�ؖh�`���O��0ލ59zLz�j�V�A�n���A���������,H!oL�cq�����H>�s�.20�_��80��k�9.�H�C<Mu��=�Xo#;:8�ѕ��~�}c;/G�cN���.���Qј6�8��\bj�in#�B��f��ܞjf��D�?�6&�c�sީ`:���ji|�RzXM�R���B6�+_49�K��|����ܪ����B�ϛ���qf�	P톇��:99���7��������܄
h����3��xíc":v	Rq0��x��f&O?���1��}r]�@�C���dCA9�>��aRY��� �cx��ѭN?��޹\J�v� ���r�kG�G�/f�ŗ�?�8C��X��/�
��ű�^���d&n��Px5�P��܄j�r���}�T;�@��6�
�or�`�k��r�����-�='��ѥ(�_�-�?��ٟ���/�1�X�RD9Z/﷌���Z�#�t����Ĥ@���Z�l!$R�aNw8"�}�� r���ë�@�;����~��E��b��K@�WV�vx��.Ǧ�cq��U�:���{k4^%��8L������ŪX�X�A�R��V,��o5-¿ݚ��ʉ���Яَ�[��c��{���������$�V�*/�@{��7�����\I�\��6�M����&�&*��~��x�sM1����Ҋ���z
�!k��A0l���\�����N�@�ne�|�ש ɵ����\[�5�o���>}gP�5�����'(cńʊ�v]N"��8�|��5���i��L�� ��$D�y}$#���ZNsy2-7d���x�0��]�HI�ɒ1���:uֿ<8�mn����D~km�`���x�U4*���j]1�[6�>?��
*F��w�uМ-֏��2�u<���ǟB���;t� �`�o>��@W>q�E�??.h�*{�I�`K2��=�^ j5pGX�w�3�r���m��y��[Z�h��]�R��<M�e�����i\���#�����kX��n�h';�uѨ�55���lr�7K8�>8����HIr5�!�1yDj-�ũ�ɨ�s��#�J�F%��3�2Rpb>'�����MK� )e$;�,�Ch�c�$�l�dҷa�q����-��j��a���X�R�hq�R
(����
�%��;)�.A���<�|����}��JV +�����~��g��h�.�)�*�a�F靨�' ��a%I���ۅ�̶k9Eh�6"Y͠�w2+��7#����l��ܺg/fѣ�I��?y�&�
�ڗ w�d���m�R,
�Γۆw�%&���r]��j��u�����IOx�ה]��gU�#j:?��5�6 ~��UL ��#fa>�v***�GG��99��[���v���4�ڪ_]�U���p� �)FMM�ɍ���_^-//jDM��N��
ْ�ݎȝ�����9<30�ZS��w������\��ƅ¤�P�?�����° �|���?t|;A�����[�u�IH3N��GݤU�f%)J�������1G�~�W�'��nF4X�?��Wp��P	.���z����2~�|��^A�I��;- �;��B��Y���!,���?t���L}�A�����:�6�X�� w����r��Ĵ#��}/[��[��1��9���"Ƈ���$J�r[9�j�?HL�Ĉg9o�E���
��׳��MMM)ǌ��c��e
y��e�ۗ�"�)�!��vWQr%��U5�TA �"��d�_Z���߄�#T &�N~�����w����d��q������+ǂC�Z;�t�r�&�@��O���f�f����ܟ}I��~좄�f�.U�A�3|������௓�4aG�8e4u��u0F�y}���@�!d�zf�R�#t�DA�ߵ��<yA���q?Gȏ���+m�#{.z%qE��)h���?�������K��	���������������_'vwv���a���G�!�|
�m���_$sŐEe�����w�=�nי23��t��3�i:���[������L�ʄ�v�^�K�G���K�7+�I!t:�r��B����.ȉ��K$anm2��B�
�����ޞ��+��`q�iK�,�B�_dk��&d��K��]Z9=]k�Iȳ2_��MO"�A+�˹ڸ�[��J�t�SP���Xʤ=��t��`"��-��O�ko��m8��xɂ����m��N����ȇ�0sY���Q"���>.6�\sb�>�'���	�obbb��*�%"Z���O��D
R1�>����<Ij�ˢL�!�}�W�����K~s���Ge~�RK�=���񪠅�$6��'?-[�m[ϥq
ZN��Å���P�^+��߹ ��"��0����}��'R����WƠݙ�fV��e�œ��5W]�T��af�9$�jٿ����H+��Ky����=�3����O��� 7���dI��v?~E�U�����������9�<Lv	b��%��.�cr��vӧ{�ϠL�Ja�c(�C�<^���,ٙ��ʈ���M�/��e��K
ɦ+Z�����6M9������i/B6O?O�b��&	`�7�.07�z�s�jX�iFt	�+;H����ze�6@)�e�|~�+����`"Zj��K��Xֻ�*Q~ֿ��d��6Ų�<Ry�n�v��j��$���V�g0˰�ˮq����)��-���]7�?+�D<B��7ji����`��('��8O��J!w�>_� ��>�[��3+*I"Γũ��G�r��b��+ھ�xllBX�|�̒�$�(�S��Ȉ^K2p�I���%J(��0��)t���ซ��y�x��!�o��R�~5U��G��������=�J�Jx� S�������4��4T���k���#۟G��wԏ4p�i���-t]�}�=Q��/:��s�W�~���w��&�K��w��(q<�?��Ix�����xd�fR���9C�A*o d�2r����xJ��q�q�拱	UmIV�v#����Y�d�J���W.�e%%����D�?:N3�KQ�+8������~��?���q���z��Q  ��u7�Z�G1h &�n�Kv�`�5���(��͑���Ռ��f���,3]ߏ	|��T�)�dy�{E�̀�Q�2;dj4�SRt���$���nݳf�Hg��=]�|N��,�|�(��/& ���e�ѧ��E���x�pD��%�I��E�'anMg$��M�����?4уCoT���9T�_�Y�hW�%''��b>y�Jo󝹺8���T�yꋐ7�"/¿ýy�}���a���dp��\����ړP�X>�/z��d�����6W(�n;�Tj�\����K���l��%_SI~���p�+��+����ǖ��d���G�O♡R�$�eN]V�:��MMNX����}s�;�y>��'2t���C'�9����B��B[�XlHF&��U�;G����Ԥ��$�)��x�q�u�">6L���K�o�����L�gZ/;#����_l��>������V�U6O����R��P�0��҇�+0��l�+�����/�x��DL��7���56��kc�@Z�_��R|�m��u{�!���d�-��?U䯹�t�P)�ʏRex5���8B��/�$�Y���Ϝ_���X%�w�2��VtA�V�l�LLzG3'&&�h�l�?%�%p�l=�!y��)�(w��4���W�.uİ��w�7��1į���MŇk[q����ٚ�
馼�Ǧ�a�!^�����??�E%pvmI��#�J5��Z��?"���2��E����,�#��#>�Up����?��*��H쯙 *����Wci���e��h���?�ɐ��7j6�q�#�+G�OJ������{�f�������ܑ=�H��~1�p!��v�xj�����oh,��D�U����m�s��Ǩ��Zw���j���7Wx�I!1��Wk_�I|�e̱w�9���
FD0�߰s���R�������X}�+����;�}�!|��O�ȋ���]��%_�@���ɬ���2t����FP�*�����S�j��8���-�UWY�:#������t��ZJ�x�I�k;,����[���ѯ߳��Q�̰dďP� kaOC��ߌn{����D���;b����Ӎ��J�/�Ԯ�N��v�KQ���ފ�����M���R^����}��(D�T��]���ӯO�s���<�������ȨX{�p�g��LTE:��|l�'���]��� ��?�ʽ�,��|���cJ�J���'%�eJS2P��+l\.n��S�_EJy�s�d���D�����F������kѣ�w�1��_���:��裸ގ�D<�����������{8;�ғ:=.q��
�����/�ww��ś�;ffPc�9.v���pL��wW(WJq��PE��$~�������ɏ������⍢F1���9��Vj�J�dh�%�\�
��`�����g�eا�������_���������ǥ��s�T|��,�k3]ӘN����+�\t��X����\&���Ӌ���h>-�2����XҒ��^/)�M��cdq�5[���/䐀Bb �֯��W�H{�.�m����z5�1��ٕ�kI��������� exVm8�f���eYF*�R%mJ���T�5��ӷ(��rZ����E��D�����D�D�F�p�y=v��g����9�j�y�pg�����:����1t�u�Z����;����v��;s�ʮ�F[*�Qm����o��~ƳH����S� ��f����c�����>�b��
�[ڔ�)�%������BV.��j�K�cA�O7�(�f{Okr6~S�D���
��w�h&����7��p�Z|d22�R�:�i����i�l����u�{y�P��R-�W8ۿ�Ѕ�G�:������%�5�,of�T$�A�}��1/�/�ٗ4
�J���{���0�f_?��O�_�s_:PX��`f�C���L�|��Ox����AP9���:L��V�ڍ����˅*�bJ�i�&�Q�~Z���E_S��.�|������?�f�k���L�]EmIߟ�K���v��!M���?R���j2s���N2f��l=�~�v�ID�Y�|�w���/Ś�����j�n��W��>#�p{�f�j9�>	�q�U���	 g!S�u����g��+�6���l�,	+���ɟ�Y�<ٰ�����@8:l�O����<;6*v�x�U7�Be��N��?h�[�]p�
]Є>8g��8�W �bu�?N�B�B���s�Y{��J�1�e��,�8���c7�<_��5�������X���bfj:���xB	O̟L�@X��K8Oݍzߊʪ����u����ӐVs��u�x03�g�'��
I�������qti���n���sȽ ��0�i��ך��w8N-��M;��"t~M�p1� :w�A�Yv�p�\o�A��:{��Xx��f�"��3�R��H9�K���>-G$k�^/�{��=lS
+ϯ�]O�,k1�͵���:e�I�9+�����G\����8
WX�Z��?<�_$ץ��tB��ѯi��
�|9\� d1�5|i;4(�ؽ�w��7��q!�Y�l�R����:*����Ԗ�^�8�]�ǐU�O��g�e]V��ŕ�I�\푨g��"��d���K��z�뜙+�uo+�ZD]��&f���� (o�Z�mE��C6��l�x+�w����x6�'�#��9e�S^�{:����i�)���?{-x1U�h��X���3��N���;F*3���#���i>x|cP��eH����X�C�~�T���wA��)���94�Ҟ�o�YB[S���),zR�+�l�6F�� ��:�S��(�MK:��}������a�)%��ɲ[H��d���a������Fۂ;a�v��v�o�u�d]�����.3St��=�&yI�7��*4&�
��x�h��� gtT��[ۤ�$�˨��4���l("���a���.��D�"e��H�e]�0��t��%0����`eR�ͱ��x.u���i�v�x���[��@%^l�{ӫ���Y�����78b����6�ȹx)\$/s�Q��K�{L�vk!��+I0�����[\�#0�.������F��Ow�#�ƭ��*���
P�hq��	y�<߁a���k���V{/d���4���[���<s& ��G�/_��g�i����t��6+����H_�Z;EB��X7�$GZɸa$ƯE�
�g�f�G5��� 
�@fg�m��x�OA=�WЦ���}U-�0�������VԻ���5���p�э�Gؘkŋ��(����p#�J5� 7_�n���G�0�p�Ҵ`��l�j��w��b��`j�������.�q�3R�m�1�e�6������_���Ѻ*��2#�Z��K�2�����/�dw1XH�_��#63�W[YW� @�r,�(��X�>���e�t��B��4��_�l?����ے��V���U��QO�NͶ!��`k�˫������ρ�IgX6d#P��sBOc�����;���oh�tK�[�Ǖle�=�*׵&�w�C1^{���߅�༴�b�,Z�ꤸ�$�I��F��.��ժF���z��B-�ʜm����Zrq�WO��U�~7�y��|C���)KC�|�IN.x>�g���%�.V��)8u �c���_b�GZ����I��K�����Qϯ�Y�rˎd���E@R�!�}�&���ҷ�X�O���� +n���h�z{�͔ۖ�M����Ó�\��鬹r�M�����R�C��ӎ5��������n���?�{�;4��{��{a�Z�H�Wy"�DB_�����a ��:���X/�w7�;�/V�)ir}S���%�o��@q�_�TRa�9{"{$�}��7կ�:����v�KP�U+	�/W~�۸2�����S�!�d]�%L�)�V�������ziO:��T�����_c~��O$�4��5nS�3�����G_8p�Z��:�}���S�M:��L���i��z���xm�p�(�m�*8�2��ؘ�~ř��hC.ģ�j�m��t�a��ȑ��R�F�Ċ!�[�|�3�%���^V����K��ỳ���2
I.8����(2a�Ʒ��/�>
e�r�Y��0�)qc�`3?GFdݿ�j� ��O�h:��Ct_�ݍ_��H�%��F�(9�1]�8��,#��o��#���������֝�D��U�	���x�v��e����^��yz�HY\�Ǫ�&���x�:/����}m]�+ao��A�l�ܹ�P��h�C�n��"�i	X,�h.�N>�5=[h���d��&��*��\n�.��� xnav�WH��Q��pB<�8v�:����)��������bTb_s����\�#�������r��k5�Oy�H�1::z��͗K�M_�[�$�Ǜ�ޏ�۞&���&����W��w�ħ7m�8c*���#R�W�#�qEڨ
H��~9�I� ���F�믢||�cc�h��o�v&�p�ga8cX��h�]��]|��7���(���Vis��Y�C8��c;iJ>��t)��~���X�tr��-���a���H��qu9Ř��&�>���Q1��P����<�C��f=�ר��7E�<@����e��f�%=�������w�$�uHuг%�-KZ8�V�ڼ�٨�Ժa�9}����pBc_:�V�b�_E��řP [2ߢ��^]ɵ�?�{	���Io_����R��|�=:�`	�b���V)J�w�m���}(x�����A��pNľ��IgqF��-�'��'wo^.w�L����57�S�	蘩���p����r�o��u��y�"�@m��c�����3&��-���^���O�C8�M��"H� )�V�Nϝ��Ȃ�AҀ�ߺ�{�r��A8
�,��K�#չd4"�:"��|w[M����p�́X���iL7 ?�tL���h�}�?��Կ'� j�;�-��s�y���MbL��	�ʟ�F2�Z��G��������i��N\�������N�T׷�օ�3h��uG�a	�~,ܦt7>5e�li����������A�7y�n��l���E��ӨW`m��ݝ�u�S�Ɔ����_$�W4�v���)Y�*sU]��Z���.�A		S��	JS>� �]G��s�Io��}+���H�`��C��~�)����kO�����-�J���3��r��ſ%da{�\�_��`ǭ7�Bg��%EN����u�d�ӋmLկ�.7����wA.u+��@�۴�3O���{x:��Xo�@Ke�2j��l�W�pQ-Q�SRS�Б��G�p�͂^[/����U�Y&R�;8T��L%����=	s	Q�ꖮ�^3h��cھ��5�X]�u�Y�6��(��Of}��3Tpg�Z�4e�M�>:!���ܤ+w�G=�����$�+��I�|�y��]&��/1E��%k��?+V��_NJ�i{����ٻ\�hmr,��Y�]�D��	P����� �H��pv�S���ٞ`����J�i0��e���Lt\���1Q��N'~�'��Xh�fdL��6�a�Ok/��)=V���j[��F ��|>��X��cu:BM���<�6$�_D�4�?/j�wk�ujHWR��H�'��U��D��%�>A3��t=��`N�1I�y>y^T�b15=����Ny�E:�Hz����D��W��t|`��A5<�NT#�s_}y��JGm��}�#�q��L��q6��g7,�ŀ��P�!�Ke�	�BǤ��*+i�<���֭�}qm��=ҝ�>W���2��9p�j��̑��Q`B@_r��P�����˃Y�}>-)2iK�����
Wj>oh6a�)��*?.I�2���
�g�AǏ�j+�5mG�A�.4��u���T�y��m�DF�ʆ�����,�{[�V��[#W�=���cb�&��u�
৊g]}�6��������J��6��{��p6C>6������q;���f�Re=�`{;��� |f��Վ �EK�,���*�E�������������������]�b"��c;���4���7��DQn`���ya�!,���UH~��߆��hi�c+��4z	� ^8_ꢇ��B}yޯbJ*~W�ϼI��L�~���X��Y�&�tйD��z���{}����|�}P�\�ߗ`n�� ����AJ�1����x�6S��L$xBǰN���ɑN�75�1�<R��ӯ�{I�O��Nv��Jg���E߽���<���n�l&h}���|J��O)�J[��}�0J������P�e���.&�AL7�<3.L>jťo�o�i���Ȁz�l��`\���C�c����,50V�n��ho1�s��鱵xje�T��W�L���zH�89ق����)oR\�ߵ���)E�IcH��~�2Nȅ��J�:+�H��(V�R�zj��p�k_Rw~�"���j�J���.w���=�V��>������ᯮ*�b+,��ɑ�i�g�"�}C��ͭ�W�'!Zh��n2��{V��:4<TDAo�@DB�����VV���VFFF2���eˀk����0�K�_�÷����{����Ӧ�}i���rëj�}h�T붣��%�y����1$�r)�F��Ɍ@o%�� �J!��{�?jK+�WP����X �2���ʔ���CZO&D�+笚T��2�7A����"�\�0T+rWw�|>�^?e�.)T����?�e�R���{+<��|�q%��V��,��{^�I�W���j4u��)f�ɟ�5hɎ���1��5]���K۟���ݴn޷����7����{KI�zV�&CI%ns r�{"7@�^���	\�e���-IF�MahW��zidz^K
:�7-�����#��YH,f��"04���7�!��N3ڮ{�+��V��W5���HoLzk����-�3�{�
����`>~������4!o�"ϻ���˗�ld+a�	!�z����_<<�CCOh׶	0���*���+�D��9W��[y��ڌb��(JA_��O�A�1��d���ہ*�x��+��wM�\���c�ʏ��" ��x����IZ���Y�-��eI��3%73eB���j��h��;�Kܐ	�K�����oI=��TT���Bhhh�$�6v����!B�������:$�^���1�9����Xrj�-�������q�e�tL��1:�r̩�� :�Q��dL_�
[�!-̽����t�O�M�i�����k+�3��]3�Ob���n{�sѝ�?���lΊ�<7W4==M��������p����;-�ׂm�)��W$�x�����P��8�/E��������f��\kn T�v��!%i$z��s��}��6�"�[u��&�y���w���L�s��5g���6����T��n���I�$U]�oO�.�X����9K��Ib1o	��:$���T���׼6Z>��9S/����W��:H�똽�x�V�:�a�6�p�5�7�s�-��?>}"�_E�{fk�����)МK�ݔ���������������JMi]���Ɔ�n�ۺ��e��8=��S���_���a��^4&�.��Zs/0Й�5���ק
��N�����xH�C�y�KE����N�e˹�~��Ԍ��p+=�;%�n22���D��+� �y�%E�[����o����- #�>i��T�q��=��ijj��G��(yz6E|/+q��ޱ�+A��Y������N&�Y�)Ȧ7��dK�< ��^�vͤ�_dz�R��W2v����;�R��.��H�?������>g����2?^n�+�0�}��Y����he]邢���#��m�hMLB2i	n�Y(�l����9edf$�5<��\.�l[v��7�u9���Z!�G�_�I�H�0s1�0U��)�<j�p]���,�l�ϧ���鯬��}S�s��}�te9�i�g�f�pr�G�c�5P*A���U��"��������^��#��MU�{�<��[9�ۿ��dG�p�j�(u3J�iE����BC&}[5���,T7����,�+�'���0��<��@��2�p'`�*�s.AC�l��=�O�&4X)��gU���-��G{���$��[<Q���eww,'��`���5�_6�//:::�����c�fO�+3��~� �7�VZck�ſ�R4�\w���?���K��=оs��.�_x�F��Em/40b8Bvw�#�L�QD�nA�����z`�<%5]�Z�AlX�t�t,����O7R��
���n�,���yHt\���� ���(�H�$��=(M���*ם$h+R*���B�ɽ�q8	����Rm9Ü<%��H0Zݵ�i�mf����B�V.C����e?aN�y��R�j4Vߙ�4O��(h�L�o7ὥܴ���m��x���#��	��^�IR�ڽ(�2�ϬW��� J����[�qq�Ȗ�i	%�^�ב:��s9�����v",m�gx�u�L�/��D��ͦ>]ΪK��ٴ��|OP��XT�&2	T�:#6,:�Y�LI\�3�:OTED[/�9nG;_���l�⍬�.)}k��Z�GG6��X���D��P�,Q6E��Z��Mx\���Q��_i,}Z�p��vϗ�Q"耎Zl�y���V��ft�ydFI5eib����(���`���WTSK��ϟ\Z*s�6��h�L·s������]����AwEH��$ŕ��?��P���c��PH��p�j�)�\���è;{�h��A�� �Ǽ������@!ō���vx�IT��Q;Վ�~w<r�#����W���û~-Vl���8|<.G��9����z�y��b����F��3/,Ę'�^TT`���8��i�r-�,X�����/qqqA���~I&F��k�2s�<S���o��t S��f�["�8H����Ff�_�0��ϖA�y����jm���@�����:�^Bި��h�Ȩ��<1~�#eiii1|��CC�vv򈈈���悯��N�Mj�-Ǌ���w`���2_�������+��,?Y� 7;� ��4���ڴ����fN�}q�f�(N�a�^�$�h�5�8V���;���@M�@�0=x������vha��ʜ?���a���nj|<{���`4K���yB�{ ���������f@�T$�h��Ƿm��p��>C��i�/2cɡ������2��Ɣ��5�S��7a�>��K��l�{��E:E\���?~��@G�K��ztUDC=�b�! P:Q WRP 111!���Kۿ̒1G��s��������1��i�4gГw�3�,k��`�i���
��$B��۔CD���{��b�#*���^ܜ����k��~�±ܨY[3�FAl�kk����M`9a�k������A<�Oj�V	���ɼ��7Sr~2�!fn82�--�����3|T���������C��Ξ��!V�9z&�	2�ye&��8L��C���n��ܿ�Y~2I��Ï���Q��'y--�%l!SW�Wa٪0g�N0t�����kɿ�,�ȸ3�lk�lg�&1����Kʙd�Msf<e?�u��oH�ȅ�.����|�+=gc��L����Ձ(�2�n��,�@g����t_v@c٨���C���H�;�����Ш�ul!�ѣ˵�ъ>���hii��uut��tr�?��Z�YK���bd���t7��:���xU�iP��3�R6��[�j,^z�jI�^I�6T�ޡ�\�劢`ab>��
�>���p�ne�M�I��.���<���{vS"L��k�/B��-����n�H�|K�8GƋt��Z�z�����`��KT�*������0Z�6&����T�\U�%��[�\N~���P��B�wf�f��N��h��Eĺ�_�ʡ��c�Y�?*@
E�p�7�L��X��?�X�%$^�p�h���*�{��$�KF��L�*�Y�s�"�.��E����������z����?��� ΍�{�=�6Նt���x���p�6�Y�y�a���4��҄Y~�g� �^ [h�v�*W���`M�%W��P$�1��c9��-L�)��$48^�̟J��3V��J�t>���ꬽ�0�1iJ�QgM��j2�����񼎆(-�ƿ����.�H311�Y���;PQ�&Fk��n׎鄗�n�y�ު:��pW,Z&��DA�ǘ3m�����<R����&	U
9��{vٌfKv�Y�~z��� 
]VR��9eA��}��)f�Y��~l��,�t�4奋�ʊ��w�j���i�Y���[3Ȣ�N�w��}��{*�
�c�V�z���S&a�/�*��wB�K�0'KE��}�GM`�P+�"�������An /VZ�%����
�����cY�&���Կ��*�m�:�!5�:�u*��n-�"2a������4�+R��D�<4��ɿ0����/{~���{3��"|��X�p��پ�&��0H>.G6߲o>���}�F&4�֒��S��8^l���z���YDQ�e����W��v*�|���Yk��#O�+��%Vp�Ǿj��ݢ��r���K�o�wyYk)�+�b���f�+���A�M֓�����m��jGfM-�\T�z|È��f���o[�~��x�sfi���b"R@d�OM*�WϞ�,#�L0�n����N���k-�\�~��F��h�{�l�bH��{���TD��A�1�Bd��A���M�������I�5_�X���1o�z,�T�C�6�����ٺ��:)��y�hg��R�E�nA��®PaY4ppY��^k��BJ*���/vV���3A�,�������S�YN\Tk�F�h7��V�N8E� ���Ɋ��NI���4ҘOC��Ŋ��i��)|�����^�n���]�X��	�&a�3ꇽ	��AV3�6
����N� ��=x=���u��"�[��<���~���d��~�FO qb�h_"���6�^��֦8��z�)��N�yWy��KǌNb�Z�n���K4rf�$�9:6�G�XXEQ�<W�Ѭ⽄s�L{e:\��?�������1���$�"��[�Ͱ��~xm��%��yg�R��8Ln�Rk0M�k'��b����r�F,���8��0d����qv�ˏ�ʦ��ת	����~��x��ͅ�LA���� �����C��7vJ�G�������8�u���L��Z=%�2㹿To>� �p�*S�NM�ǖ1뷥��D�+j�Et\��QcUae⎛���xA<��TҶ���N�;�Q���~S�ma)B�����ʽ����/s]v��W,�͖����c���t,�d��l�H��8�W����	���[3�hK�/U2�����v蝤�h��n� e����#�K��@Ơ #���ji$�ō�06U�D3�L;�,�������S�fx*���0�B�;M�f�����g|lS}ތ��E:�g���O|��1�R���c�2fZ6��K#m�� I^_��T�2</��nyhU��l$�%����fYtj�&�tb�a��=���P��yf�����6GX��a3z����ؙ���o$��Nj��~'��!D���m��\��|rf�y]��o�J���I��r��T�*�N�(��F蒊��0�Ն*����aj����h
~�B�H�MM�lbu~wDv���OI6��Z.+��w�>� p<%�a�s��]lSӓ������8��J��*��$��J�5�Y:�k;�����|wb]��<�@\��ւ����Q!����x��6-�ZMoĊ�����+�c���y+��H�A� k$I6jcP���+�cR�cғ�>*9 ���kS���+�> �(�ZI0d�������Ed;�g����L|�)*�A���G~�7HSr��!�d�a4��2���a���LD��bW�#�Ἳ�����z�����pJ��
ѢK����[�,C��-qR��W=�>�lD�rv��)	DU|��X�M������ի6O�B�A���K-�5��<^^e�B*/������#o�Ȟ�M؜��>dO�e��֞�����D$��""��ͫDS���%}���K#�k��j^h��I�����޷�tF�3�6�"��������u�':|_&V?^j�{A��b���q$�m-1)��:g	P��SU*��n�֌2Ǔ_&09��&Sظ��Y�}���zk�g�r4�:���?���)Z9�cA����,�n�ϹY�@8\_k{۠�ZmQM���=�N*�>��Hp��n��
s����j� <)þ,����j�Y4Js/�;RFM�B����So�R�)ZI|��4�N���Oz
����Z�F򹟧�ƟN��B��-~S��֏\���X���9���*�4��h��'��˒�7]�1WTD����-�9~��8���i�㩰aDk%�t+�r�z�X��/�Q�F[I�V�s�o��(/��Ӡ_���x5�K��Z�.z/���Es�_'�W��Z�P����"I�=�~�Y��o�Z}�*�e��P�v�O���s�*�*�g§�����OP�h��t��z�g�	�C�B��l&���	�	�+��h�/��N$���/j@.�#��=S�u��J���������Jj�q�o��ES�9�����;#Ֆբ�>�H������r0��w�:d!SX�a�4���H&� Vd�H�7_E��p"{K�Y��_�[�Cs����5jO�^2�DZ��d��|�z+I��%$a��̗)�h�9�r1��$�Ht��y�]o{rCPs��14�~$�-1�^��~�>���*��Y�~ų%�<a>���ר�{Oj
.&�����xƍ&�8����(g,�?&H��;�k��I���7&��-��u*��F��\���:D�����D��PC �P���pq��|s�˂����&���������n�播^�LEB5Ԟ�@j���;�Ԭ���343۽�,��`xQ���Z���A���t�q�nD81zjQj\p���A����U@���Grg`v���<Bf��4̼�;�Ĵ��3g�C�$(тxO�#��o�l׾����ֳ��������Z�H�Z~�y�v[`C ��z�u�	F���ms��5Qaȍ� �z\ ϶����� �#O�0}����<=��:3����Z������T_�V�0�J��;����pp�n�2zl��j[~�vs�+�s�̂��A�缪�Z��߱L+��{��Y�����=,Nb�Y
Jz�&ۡ�5�.I���b�M׳���[�5M}n�m=��߈n)�dM9��?.q[�9[H^3M1�h�K9��*�s�b��6���5�i��BL��n�~��S�."� R,�g�#Sׇ������� a&�c�/�M�{[��Ҡ ��ط��#�VЭ�qج+hA������0�S�����4F�_�0]�\x�=%�߸0>�ս���(Xf;c?H\�ءp��������g���B�dD�dd�.(��b�o�|�k�G�J�!HX!�!�o��ȃ~W&��3n>FЂ���`�WP(��P�r��Y�m[�rѢ���p����e_�H��*)+��>���1�"�Ԗ�Z�����F��Ř��߳[-�Ө5s��i������m��?�E�#w[={�o;=�(SB^�YK���xʍ�hRkY�OGT��
����`��H���L	A ]XL�dho�Iz�j�z���27Z���eu�}�(Wd	��L��.�3�k�V^�Ul]q��wQ-�������ᶨ�	<볳eVA��W���%L`���9�����`�a����W�9�.HN�V^��k��N �d�x�j`vZʎ�$J7i+�F֘7�'����?�0�����X�2fm�lz�D�AUh����<Q�o$k"`�J���*2� z�L�k�4������FcUx�.��,�V�nw:[-�u��ԁ�(4� V���|�a���L���i����}n�#�hI���<@ADZ�LQ.d�ꙟ�"df*Uz�#�s��.�O6�/lL��3qW7jK�1F�ԑ*����{�-��k��1�JqzR/����ZA��]���]�����e���+�7VvM��<��G���+d	�|1����<ޭ�J�KJ;���3c���D~黸������ƿ>�Q,_�S�?�ROpfm����1���$�4�aM�؊g]������8��wy[��5榙ػи����@h\9�+f�+ �B�Є>��Ou� �]��X��4B�>�5��p��0x!��8#���U�Xm�r��Sӌa;����O�o���~��QB��[�� iD5�`K�Ք˿%�h���+���nܻ�e�JԿa0�G�k����`4�`��W�$'����wu��������~ѠM^
���l(7I��9����b�����+�"��U��B?��.*�U��F2C'+_���^S�!������K��x{4�����^wx���r�p�K�&�{�R���gN��yPIa�+;�j�16	��&x�W�k$4OO�8����ﾍ�Lb�~���҂��]�Lc��b�2ZK�D��:�.�.�V�
�L�#������)L#�����W3���E.,\x����x��ׁ/����i����OL�m�������=O;�WY8^ljyvЂK-K���I�@������0���r�_���42��v��.���QQNW�J�n���{c�(S��a�zH���3��y(~�6�|~��`�ޛWV�)��c�G���.s�����(8�W��s��Yޕ�^��a/�ø�i��MFfM��Y�r����꣡J�x�m�"�]�A#��`6��)dB���&Yƪa%�H3>��}Y)������3mZ��v��4��0�ǘ��N����u]�{����y���{>�{�}�y������.�T��((�}���7Q��;�����uJ��럅��s��*��Ƿ�����7���������rT�� F�2�@sT �T «A4���Bv�0Y��ԡ���7��n�2����J��dd+�7�(��sV쳇�ǆyU3+�}	��Oh%Zg�T�	0�.Lx�LC����󤇩Vq2��GkV�@�����A�S\��u����ss��$��9?��{x��.$��MC����3Pl�Ԇ��_߰[zЩ��U*%�ͣ!�����l��9��Z9̝Ōw��N�kȝn��M_��DZ�)�P���j�C�"�ӅB���Z�8}@u�vҙ���\I�z���jd��989�ک��㝘�ؿn��æ�E���:�D�s�ł�W�g�D�N�c��sן�U���=�\g���qٓ-���Sh$ϖ�u
�"u�})	6Z���$2��!C����w6LI�|K�$����';�2�������[B;k��u�j�1@d-�����<�>3 �2�t���\�M9�o�~�ǔ�ax}�������
�.�����4Vʯ�*l���ǥՀ��o+3���S��T$Q���]���,y�K� �<[~�s��hKU<�}��3���T�0���>w_�{���Lc:��޴s�G�3�o�u�+7���"�T�W9)���Q��\�"P��c3e�%�kXx?�1)�3q�wqq��?�EAI��{D���8��>�tR�*k
�����CO�h!N񨯜�N��0�����pe��*2��f/X0Rs�W�gB�yc�!��`���#�=�Wm��\�B���7kBf��U�ۀ�'EȌ�5��cq�R!�ށ��Q��L���x��v�xPD1sy2��dIȧ�e�]��.��E^���8�NK*6o��m|#���0� ��rh�M��B�n�U<��+@�	�s�R�\5��{W�4�hpp�_44䠖�h\fb�p���Q٩-��Tę�9��Ֆ�&i�hݏP�}t�эN\j����n���4�dT��!�#q�ܔLz:�nڢ��;�͊�O4�H.D��v� ��q��D����AY��B�����
֞J; =��l�q#��ɠ�k��H���聶�n����*�׻$?�-j*?�4(Z�@���@�ȶ��u��v�S0Ns&�e���a.����r�%x�ꉴ���ڭ|잇	��zxL���)�]���@�!��E��i���H�]��L�G;���[�`��lsD{��|ɮj�z)s�5�̈��m���K����]uٙ�hk����2,�тԮ�;k}��~f��T��i�Z�"�.�]ǻ_�z����Sr,�p	�⛆��b�;�����r%�G�ℵyG����ê���Q<+[�l��Y\"�e �afr���J����S��{ &Jy9k��QUR��M%�2+ѭ�206k���9?�J{�B�p���t	=�/PK   ��dXWC��)�  � /   images/093f54e3-331f-4155-80d0-fca9fbcaa25c.png��	8���?>ҡ�)�T�9�TBC�,5��A�(Kd��/�q��2r�fP1ɞ�0�Q�
���=�k�}��~�z���������{����y��{�_���ǣkښ<?���\�����.��~r��>9��"�؉���]���u���K7�0ؑw�v7����0�='k��-�;0��v��h�[�wN;��ď�?��
����O�h�O� ݯ{~bz9a�.n���(��@�n�OoF�������_��v,ȋp�qW,��!��U�Է��N_�W��+��ޫ�}���.}�s�����}2lTSr��i�� C�s���sJJ��i%������鮋��?�������� T�źȜǾ�'w��A�t�+��OhEz8Ϥ�/e�>���e�%���%O��'�3W�L�����TV^&�o^����{��b0���.+Ű	�~�8�O�m���z�K��n��矌�t��d�D��`���JJJ�a��8�]\o7��N���;�Y��Kxrt�
Q����G��jm$M�KBS�='{�VVX+���i6=�˯�hT��_�1g���a��p�ݥ���6zC�*��4?,V����U�\p�{�3xc�w
C���\�"��	Z6�{��O$�O�(����Wj%�X����K���}�u�=���'�5�^%U_��~��!a�@G����1���̦a�w��W���4�8�$,䄞/���v�G�����^�-^CY�	�S�	�n���!T�17�!~,){$'L#Y'I�c�*1��9H	���|$��~��P�M�P�?%ͬLZ����{�OY�'L�oUۿH�H��������e%���OƯ���CkBW���Ou����Ƥ�n=`���C�\������Ŕ����ORŖ� ���۟��(����򣂒WP0;��e�*m>���G]�
�i�jl喨4eX���[\Hk��������6��ņ�\�B�m;�=��U�C�89ݻW���sv�~7%�f�J������n�2�oQ����u���^ۗ��% �5��£9�Z��;��� �1����p�`�g��7�Zt��nf��J/���DvE�.�5�b�`=ۥ��"֛�����K��ͫ��C��zCq'�sN�z�N�����j&ӟ�Fs�/��!�;�p�ԓ��8�L�aOǆ�{�����BT�}��dPTbߘ{1�K� ]���`��8�6JqSV�K�O���0�`u'��oB-¼�E��a��+��G���s�.��/�2��|cB��6]�`�2{��TW��wAR>ڦ�ªIϕ�s��}�z+/��Ra@�;�b�.NӍ�;n�`y�O�X���V-M����������D8`y��<�D�Z�5����`ҵ[���X8>�Q�+�Y�m�L�Cp5~"�i!����a�
���	�MO�����B�"��2�T7����\A�I�o�}8�àq�`_�K��w�.N��<�_��r+���>�m�0!��	�?���c]dkjd�9�f};OA���HGX��[[�klHR���B�I��N�-%=]�$X�v"ɑ4n�<���v�{Ы����1�����m��(�_?�'t_'s��n7�Z$qR-g�}�����
�3�U�	�ۉ�Bk��c�4Ƕa��?��d'L�_�� L'@\���P�>���u�y�f�O��1;arQ�	$|I�KՎ��^nKɳ�4X�,D�|��"93��"���$�7Y��y�������@�N�K�d�ct���}u-�D��g�w35_��e� �2ty���dM��E�Uಷ�'�;6>���X/�I��>�ѱ�*&��7_�~7$c[F�O-n"Y�'������N������-��C�*6g�uv�����'z
	��r�/@B����p�\j>l{� X��P���z8�&7/o_qq1��w�7~Gg� �5��O�|��Ijs$����md��41��=�Y���E"��ll�]��wӵ��x�aΗ�����b���w�{q��lO��5ޣL��3ZVZ*���L��6C2�\0��`�}�^,��J�t��B)��x�K��x������$zU׏׌<`ۋ��s�.���]�J��ˁ���#�9�!@'��q6���$�����/%e ��EM���ˤ�(r�1��zI"���� zZ�	�����߾=JM�>����WW�e��Y���9m[9L�(�������[��K���G---����f9�1{RYQ��&c�.E}9�]�Q���{K�r0?��%2�%�:^3�YO����?��dH�UND�k�@ �lz����S�9��Fp4�����h�]�|/�5�_DJT��'A�����^AW�H������ b^��z�����z��efeU��Z�D"��e�wI�o���Һ����%!��k�K��n�^������rs;k����W�+���Ȉʷ��o���MI���Z�]��󘻕���w�C������FF�@s�F�j��[�,�HZO+�qm�n���@_�w�{����f���w�_��6r^�@�I>pC*�ӱ���q;۞=�)�@e�A1�E#I���+k^.uK���'jM?f9� 8�� S�@�T��.��w�=��U]dnI�p���{��%���kS_���S'(,�Q	f��.�����f�kn|���Q�+#��
 ����g�T/�����Y�y:a�x�[�%���*����f�4UQ@!/�2��p����W'Xk����u��ӧ��e���[��S��7��c}:[w��1��rv6�b𾿫�a�g O^k8��<���f�\^c\�s0���Uv��w�
ܲp��V^w�� ��;��?ݨ���MC� �M:�M� C��},\K��RZ�B�&� xVZPp���X�{��E͎�Ύ���S~�=�y�tWj@�XV ���<G ���ؓ1�;Zv���5���Ά�V��l��&Z�	Jh�^��kd����o������������{珰���6�)���i�,w�&o�@�X$Pڡ�� �4���Fe�)<�8��O�!*7141	u/6U\�� +܉i.��0��O� ƺ�:w���f?^7�^,sp�f��t��lhf������8U /���@����l�T�	�5��it$�ޘ��%�O)>������Y{�h���t�����	�m�ja)P<͇]����(wY�o-yꔧ�Z���x�[�'���<��G(�mm��	��X�����Rp�[`)}�ROG�H��F�E�8�3�	]��}��m�L�Z��k}�ES]�w�hA�r�����C��ќ����.�&��-uC����|7˴{a֨��fvXq����Ps���<{�#S�Z@�S�d2����U�%V��ә������q��������^}Avֻ�s��j��A� ���f��U�(V_�N��j���3E:�SO(7�|0��5w���P\ؿ.,<�<g���� ��Fe)�X+H$���4����F_YLb2���D1�_ל��.
u�ԩH���gv/V�O*����w���AS'��EA����K�W�"i�Ts��_Zzz �XPP�'f�V�u���7��:EvQ��~��}]i�Z���{��oG�+��C�3�p��HF?v����;<=�Ez�����&[���j�����$]�A~~<N���ie."��Je���]m�=ɧ<���B��p[��k(���Z�g�_ou��Cj��Z�7�]��:�/EEhV�Y-6��L �W�u_�X��M���y��J��z�k��/-d�!B��������ۤ�3�6hBU��]��4�,��� ��%���^�B	���������6�F���ă{��lp�őhF��Øq��~�,�G	�k9-WvĢ��p�@SμL]��.�bU�T�99b���}8�u�HrDq����\��j*bcku�M#�� V��Rh ��qprR�z�"��ž�AQ��ĵj8�}}�EW�#���}l�<&�8�Q���xr�wR��`��Mӫ�
�A�M��(ƭ���M���o�������)+۞$�ƶ��J�%%E�]}SR�;j���oԦQx�])== &8�����)�J���u�rY�o	���Wy{��_�r ��Y��=�6�WC��U��<�f�i"% �k��3r�"�zC�����gC!�,�J��b�~�����������n�	�6tBHB}��z�����d;����8GRdg�w�c@��
��l�����0YeNl{JJJtqեӭ��d����(�ȧ�����tl�3�l��vd�gS��J��I3����?ͱ���6m�c
^S��IV=T���ODy��t_s�V
	�]���+�}!h͟;Iv�f�B]Gը} i���4">�)tf����<4��:��J�'e��-�([.��z��.r�)��M�o �0d����wHGܚ�/f��?�T������K���k�=�����o ���>D������C�5a�]���+y��_�������9�f��*�;ǃqX�U�^MO�p��L_�6�p��͆7S��> H���j�8}�N� �V�5���ւZ'��QH�������9����Lv{�M5���;�]:m��{X�yx6�
�U���ꦭD�X��l �@�T�D�)�]��<*la�PWo���ux�j��rF��!�Ne^p����O�̸�t����_�YC	R4���&���JJx�Y�.E�ɣ��S���p�j�T4�J���қ����g��.�Q�'���E�'�Ν;WF�삭Q�f�j���1�6���ک�<�éQ� �e$��ݟ	Z�Ys3��@%�-bz:T�)^�/��~q��SfK%�/��^6�ʯ�$�DY��� �O�5쳳�SF^Wm�+$Q��\n�$ �k��#؞������,��I�#����@+p�J�Ȭ�>����"̎'�~�����o�ċ����GX;]�z�@�~���&_֟˝F�49��Tzϒ�V�����Y��s�3�g��`,�H���k��yl�=���9>�745M����j��Ry��w�TB�M��	~�[� ;��`�h<Zg��~�v/wu�4����6Sz���J�$�ZҕђH]�t	�訥#P�>]�?K�����V�Q�;-���RampX�Ř_ާ<Q�hߤr���R��t�lΣ��D�Pܪ�=劲�|�������e�]��cl��֯�R`�,}�6]���.��Wf��\+x�+��W���s�Sk��q,���Xwi�Fc���}Y���l(��+��O$.i2P9ި��҉0r���#�h���ȁ��co�M�͡O�0)�J�[��� �������𝮟���S0x��1�a�tB9Ɛ�`�G B�KT��Z�� ����d�|I�u��]jDؿ���*@���v;�i�U�2<T�}�rjk�e��i��������Q�+Aw�&�e��=|2;�����R\Z]�:�$��@�%�1�z۸YV�(P����Ŋ��],�|M�G"*��q�j��r�J��,y�k��䐐?�#������������&Y�]^U���3�8^DO,y�w��\����>V�<߱���(�@�ƠQI�k�,�س,//����,?%��1��˫h�g����Է�S�Q:b���n�s�{�wͼ\h|�"���I��)�i��+D츷��� w�Ә�i���kÈu��u`�����$���v���-T��T,��UE�K�X�Q���g�P�A�fؙw��a2@_��5��8�'�fyՅ� �"����ay]>�H��'���$��[��
&�Z��}��*!Hu!�s�x�h(��ݾ��. h�P�s�*?��_�u��Nm�ݝ�~�C�V����������W5S���7�x�L��h��TE�|�A�����A�#���'��ݓ4[6�Uno�vB09;���L����;��q����d�I�H^�77��7o�G�z����O~Lf]g��&+�k%}pM|$��KM�'c�Ck��Z)G��B��Nii�E��ih~X��|�~v�l�r�M�����J�p�sM����bta��I*���f�����\W��,�c+$M���g���Lk���6;Zq��ɓ�c��m'&&X��o��[�VL.��dc�)-���%���w<���n:���R��l��H�cW��)�M=5��KA8�{��Lj��r���s���$�}a�֜_�  �S�O��w��>�ɂ��B��������5R�Ua0B��[�2���Qq�9�#�o߾eZBlL��o����/ �����������X����gO�?�7���_6����j����H	�xr�M¹�-g����3�ƿ1(ZӨ��i�#�X��IYQi��(�@+h�X~����pG��E��֚�(TU[�ԂH�}���S�F^��<?k�PEU"=[+~�C#,�\����RqQ�M�\�O�0�
){Z�5_������֞���V�i��mvv��	��bd^��I�ø{n�x�|��333:P�����A�p����x(ӎ�����AqmN;UO��	j?p���|`�g����� 5aW����'?p��%o�
MB��ϣ}�`FisؾȚ�7����nM�brA�
�	���/t�2¼}��Y�0a}$cIS�o��t��R�A�(�6���:��� �<J;�d�X�bB�xZ�ܜ�_�OhP���=�oI$-�p1���-��'� �"�(�U�	]����^��9hbs����ؐԶb��:%�ؖ܅?���A�TS"�n�i�'
�P76+=�-GRr��fjs�U$�~0�&��X ��KӻZ�>h �q@�=������J�λ:�A	����
b�<� ���ݹ�_[|�E�jf�)I>��� ���U�h	$?qq������\$�[�W�3!�d�&<f����Ļ!������~qm ��6|���TLX)���<��Ьw�?�-�x� �1 ��!_���C�p�r�~�M})�y8�7� ���;;;i7����h���(TPAHK?��꿇+�U:�|R�(��
>8?]'˞Kwu�12�~��Bo�m�C�O`i�;��@��:نJ�V���#1�!����>��2wfD��t���^��s���0"�Wh���[�m��W���-��!�`��gc����ŝB! ��84s�*��IQ��@��8Ȝ�995iz�� ج��\ޒ1��o``u���o�><���[�hȽ�����M�v�@Un+|��Ǟe��� l5�ѱ1���k���aY��T78VFy�����/n��R"�k߹s�#Z4�4�R���c[^t�BF�wS|�#I�n��Ѻ�)
u���T'S�6����w�0� �����/��h�>nAd������?mP�}���M���㝅�@F��&���{{���e	���Yb�����A96�	��='kYq߶נ�2��7��(|]�_��J5	�Om�����r�;G�����fF�6�]��+֘��}�H`����у������O��(t�?���̗���vh�
��2��/��
Ƚ���p�߫�NG਴CU ���{"��`������z��7\&;{(�t�u��V���D��+�n��SRI��R����n��}��V�翐�����2gA���r_:p��(� h���A�@�5T��.�4Y�St_��k�ׯ�����`	���F�s=S�a@_���ͧl�����9�k�f
�{2��Z)pڄ�"�<�ޅ>����% A�
��i�t��rmSu���QI8c0TT���w�}g�w�燼*�
��]MG�A�(�q�F��IԂv�<'��y�%l5���l���b�V_�P'�K&��!r�^��%�}�i�}�=%2���Ջ]{_dgqx�>/���TF��=���+��z��h�s�n���w
��B���u�:dt�P��x:����ms9�k!�t��Y��n���c�p��ۭ���T�is�-���R���w�@mԶ=�_V\�x#�[�-����������`�ݸg����@�b˵- a���}1v�bon[�]��_���&, �b�a�7�I �Љ��	� ����
����䓟�1j A7Q�Y���F���Q�(рN����goG//L�a��� �,�g���:8�uX��7����{9x[�?<�z�>�/~�s<�?��m���Y]�5�/L��<�ǲ��o��oT���u��������޶G�8K�6�.�f�l�W���t��Z�~���~�F�����ȝj!�FQVgdo�S�(��(���y����e�D}z�CдI��Kg�˶�I��k���/�������ہ���@���o��ÓǠ�`y���
����}y-nVm[qLbM�����A&)�9����I�������.4�՝��WĦD�BzDm���5�֗�.�k�����z�e�� Ɲ튌)(2����5�#=@���S���hZ0C�O2VO#�n���K;�T����\�r�޼��w�rq���Ѭ��e�D[�+�ڶ����qO"M�-<�}���L���]��ҷٗ�SH��^��ČG�2�	�+[��H���7���2��;���S�mn���4�͛�O �a����.<���8�~�g����gB���	�׹�N������oR����,L����O��Z�4{��/�%on���3��E��Yږ������:�z� xݼc�Ti���%���JܰR g̚@"=�o0IB�b6l�켖A� �8�z�#L<ՈY�:ѹc�aa��@\˨�V�{m���n#V��x��>���<K��au�h����d�gu�;u����8߆y^�"��@�`���T�1;wI�/Ok���B�Dܐ�����_F�z�!M.��u��K���r�%��OV�Ն�*���	^��~�sbp��&Ӊ�i�B^Se�}�q ������[���81�ǘ�DM�"�D�w��Sp���G��D��D�����)��4�T�����::2z��� �1/yN��1i���3�1��!�!�?"񗈤��}8o�5����5(1H�(��f�����K�:���r�W%��TWDۋG�(��^g��º95�dro�N�Ж
�
��D����!_语z�X~�F�p"�^�h4;z"�&52I��������F#%[ \��Ng&uY�u	3��UR������j�Cʴ����kJ���5�Zn�W���O��T\w�B~s[��r��h�&l���U0�ъ���������u=����(�W����FVrp���o��M�f�-��{_�:/�K*	��	׺�l��&C灧�������}�����*���j*�uը��ΟF��1�_0li������O��2B���U�e�St|��_�m�+��;/�N���L�X0���U{�ét�V�Kx��,|��/Q���W������NiV���)��;�TV$&X�q_gʗ��Hʝ�~���{68/'�^��������RC~���p�LnE�����bt�%���qF*Ӎ��Z�EK'�7�\<-ֻ@��ef(vu��ZYmyB�'_���Ǵ�3C�n�S�O��J�H�g�B4����,�����n��ު҉���[� �=2�&�mU��}�����_%�)��	��U�;����3�qY��d�OUg*�?:o�\S��w*9�Zx~ �q3������%��r�if�W�x��*o���R��	!���)7�/�R����Z�vJ�az��a��V���H��A�\�~��Y��vإ!<ĳ_wΡN%f�W2�>�2����P8���`��o0�'a��_3f�P�h:W�6�	�(�k�2v@5�?�4��pd�!���X�����VB�̡���&U��Eդ�(2S�?�McPi�U�2����5;|���&�-�P�њ����+�����4E\������//	o�+�Ӕ7-xj ��_B�*��f�/�;�yd"y�S���Ā������1�q�ܚ<<��Z]ɧJNm��ޯG��9�1 �I��i���U����y+���Y�j�;����307MU����#�(юYK�����vO�h�x�S!񥘘��~��WGK����>
��$���m%�JB�҅x9��f�g�%�iz���8��-���b���fi�����u˯'Ȇ�/7=�ߤG��i��؊I���6��ϴ]jiӸ�s�_�ߌ�Q+��<3���8sO��ȧ�ZR�7\���q�c��*q���sZ�����G�_O!����5~�z�Q;)w8y��Hd��O�o� ��9�S��&�v�`^�� ���q���	�#�m淪��[�>�4ɼ�(�$PwA���� &�<H���rƌK���$� ��.zJ�C�G�m�߿/�3S&�o����^Xs�>�t�k#�}V/�\n5����X�蛺4��)���+�:�6���������¢':7����蝈W&������H��ԒK�E��R������ϻ�8��\W_�;Ж?�������;��[�B�ԩ�)�Z���R#_�g(��dgg����S·"�O�i��vE���o�����!1�1 ����k�_#����{)w��-!W^J� \�#��#�EEýK��i�=��/]���xxh������i����[`糼�^�o�0�LMIe��Q���G"��ej�I�:��j�$�]ۓ���QQ9~\�i���8,6q����GDD�p@�Ѯ�Vz���сJ�c't�U�ȫ�Ȋ���ݽ�|�U�ik�x�u��]XEj����&�ʡ!���P5���p��+R���ے��(�e�Z4�@c��.���D~e�q�#պ��N��>!���n-�șH��<:�C�rr��� Ä���_�E��'�L22��<�>>>Z�� �A�a�X~�b�S~J��z�~�E��L��-��&V{�Aȧ&����Ԅ�W�����.���_��4d���zx�ė�i�ɬE$�D�듹yմ��x�z"惤
�4 =dm'Iihjj�^��L"���T���nH���{%a�T`9�O�R��7Z^u=�U�+db��C
����A��6NJ��=����)4,,J;�}�[yn�۾���p��U%^�Hq��CPV������OR$��mR����o��`���JC��-�H�u�B+F��Ç6��ꁷ=x� �,u@�L������ᝃ%�vmc����c���O%8t���������^?�����کS��[>
y�F��25���hW�ҁ�&
�^��lfC@Ǐ���W��;�|H��ڝ1Q|V?ʳ�q����9^899���Q�U��}�����2��3���v�^~(����&���j���v��ỒWJ�l���)�cv��L�>���H(.X}$w8�������`"$�B��#w@(��k>�cZw-��"k�����bm�%h]�E��)����ۿ�ل+�У��ī��-4����5I�Y��tx�+^'ܔԜ�4S%4�5
����l���U-i| �L�����ӻ��[�|0�	���c����\v���ml������3N�_��Tg�H�UY=����4E*��������i{.^FZzom�dHYY켃k�<��v*�~F8m�W�9�4���1��o%9AϿ/��z�Ds8g��,<���z���4�A*�v�!P��}A�!2�Ǥ�`)s>�7�����W/N�ʥ�:��`�5Oԇ��ntGC������^����T�������C�����R/�@�o&��k�B��7
��D�7��[�tᲄ�)䬧�|�����7^5���Q��L�ʕ+�==��TL>0Og��+5�6B����̺���3��.M�ូk��ϯe	?��9O�o�f�7��j�MҎI��sc!��ă�+���/�<9�~�5�+y�ٝO��3�[;ᮊ٘�j6��~�o����W-ws-��E� v?�[e�|���B~:�~8,��*mM2���j��Cg�(\��H?i�C�v\�+
�#���xEnX /@���-����W]Ԧ������ˊg4����?đ]��=�{+7:��z/�Fr��3�>��@m�����ſ��E�eu�9^4��l���V'��s,[i@ἆ��@������"�B��?<||��fR	2��+[���Ow �pRj��w0_�m+�vu�-+�i�2W������ye�z��g��Ď�I��KO~���a��WJ�yp��Ԩo�Y1��`��%2��Ǿߴs�=�>(�"�	���o��ci ށ;!m�.�J��e1�oAߪh��0������a)�.�}���I|`�(X��8��EO���&�0zéVׄs����gϞ�
>Ua>�g���;���VU�����M��BӃ�!D���7wj-�����9�K[Թ;�U^�	+� _�q�X�AX���\Y�mydW���o<ԏ�>�}�z�jk����-�!�6
5$�ғ�T�1�8����"��pE��Ґ�`��eW�W����ŋ]*�5Ր��iqB�T�2��=���f��iiJ���z����&#���/���[��t�8��M��h���#4����Bv1�py�85�����j�Qe�ѹ���t��FE6q��^%S#����56==���S!��M]ş�Պ)ȝ0�k�B�Wͥi��2�u�`J�篢���w�J0S0�Ƙ8]�gnT"a2vy���>�q�{u��f� 0�|Z�ݠ�k���0�R]أå����������N�i�c] �02�	o�./���q�i���ʒa��4悙J
�Sh{�b�l�Tr�5�����dIř�W]�����bk�@i��4_͵��+|�{_�bֿ�ߑ� ��jqj��[Q�K+s��AE�M,�E���Gj#\<����0���dM��ORV�bJndE[U�����<z�h�A�/@&�~B�[Va�X�>�n�mE	�����:w� ����d����:.��C�K�:t���K0�����3k*I������Q$��󱀹<���V���R٥sm_)Xl<���QU��^Ԏ�� R^�,g�[���9���,�J�YU#�b���I�dA�;k؜UDh���F����<3�<��6�;�G���n��$`F11�**��d9�%랼#��X4���f�;��86��4�IE�A�to�����k��"�4�	�E#X&S �T��鈂�j�����j��h���¹6����� ��	�B�.O�-�DpܕY淼�/�����߅�' o���h!�A�|������O����m�h����v���1�l�I�72�m�ւr��� ���A�4q�vg���/e��?@�k,�ȵӻ�����A���3Q�w�Ų��	A����3�{yL�5zE�������rT�����/Y�}>��fZ	����\bW��6ߦ��ʷݎ&˙({Ǒ�H)�>�'@|6����a��E���Ϲ�X|�AW�m`n[���;��Ż̶��|��S�Ar;�Sr�
coǼo����щ��]X����og)ͦ-�8a��O
҈ޫ��g�����|eN�K��%��ǽsg��P3uB�����V'H3uqg��&.� S������P�b��%�M(�P�#R:��m�"��j�I�<WU���d�WWpŃ�-���ϗ��r�\ANU�Gw'M֦����}�c�O w1+A�m{��ܨ�dNz��D��D;j�|�?�����$/:��4�d���������QN�ϴ���Dp�FJL̆mJ��׃~�����5�ة�RN���
����A��j�F���A�e�epϘ5�H{!����]�����"�&z!��#�1�/��ѲL����k}�F����KJ��'�K�c.,�\ ��'X��>@|�Jy-P����q��BG?���(\�j+o)��,�㥩G�LL���qI���1���t�9B�%�Js55c���V�<K�R��H�"o��E��B��zsZG �7r=P��~Y5d�eU�Ĩ���G!�i��P�J9;�7-^.	K�Vݲ���g���[=A+v����|ױ�A�7�o
K<iw����:'''@����4+%����U�h�
�n�T�?O:)��U�-�}XT�Ջ���4i�_�}�k�$M���2J���i~�KX��Ț��$Kޯ�$�H��t��+[�"��O���r�xaԾ�����M� �h�H�'�,KF}�Ň�|��kj��+F�í\oV��+���g��8��(W[9.w�^�5�Dݝ|�ar�y�}M���Fg�E��C��ے�S��.�����ch٬dNNN~@h"{�ы�؃!���e%��_++}��$`���i�J&��t���.�4���_X����vZNR�>y1�iL�!T$^w�'��S���\	u��ŉ�!ϘZtG�4b����Ȉ9�;Ӥ���Ғ�J�w� ed�y���a��9=zd2���ZZ�6KԠ�H�{#�I���T?98.)D�����J�s��sj�����{��.Ȋ�W*�.w,����/���A����B���͜Mjƃx�*M�F�4�.���냺vtl�@�'IY�B��
fw�u�neC�X�:V��wv1���쵻������G9��W=A�M��q��-F�N4��������Y�ң��VSID�)@v��}�+x��F�}��=Jfe�1�.�3��,�^�tu��#��w~R`�W�WAAA����Š�ڬ�� �R�vQ�]	T����6K�Ɉ�-T�$/��<�]�Z�ዬn��IY�?2�����!B��e����<��RDc}��0�)���볁	����>͔H�z����݈׋u������n�(T:q��C4�uh�:�CʩM�u���\��.����g��"��U�!(�����Vۣ��0u�L��Or��Ԡ����~(��E�]��>?�i_��r�k�w_����(F�.6�t����'��(k�X|�o��꣹��A/d1��b��qMh�԰�ǡ�
�\��#N_�?չCR� �E~s�2U��"wl���E�+�_��Nl{�����s(��<:���2W��l����<�rW)�8���D+V��*����Y�� ����v;!1:�0a}�؀�X�|��U{��n��k�j��XYN�p�oO�.��EZ����]�B�ռ���uv��&�3d�5��+�����\��{��*�WEn?V���d��k�8x/U��@r���>Wo��@�ӊ=!"�ǫ���o�"/��(ned���7.766�&5]6�d~X����Y�ߗ/���m���c"9o��d��"�1(�A4�= 2� "E~m����ņ2��AYM�OX!�u����Hƹ��e�Ӈ��V�q��7�1�m��W�hD�+��B�=tas	����Z+��l\D>��-#�=o���*�0jݏ�W���_�]nr#��RQbce�c���Y ���\�:�eu�ۄ���?$ٹ��?��w�Q�0K^�L,&�e���%�n&�7�&����f|X|/��I�����1�sf�x�?�v�Ӈ�m	�e����~���@�/���$���Cm�6�G3��Q5Z�n��� c���������F��V)�Ŏ��Ģ�����9��bE"���k�j&�w��cO�K�1��W�'�N�}HSUw��I��|�%z"ᬱ���_:���u$U�Å;�(V�~�Nh;l�X��Ԑ��P�F�YxΉ���S��.~��*��	Ct�8�2��s�X.j��:�^��2E:aO���R����a�T��Lw'|�"�l�i���gɵ�x��'ѣ�6��FW͜qd�F�i��������x"2�5+Wh�u���Be����I�t����9�VkjMt'��V�`�(�@ݻ��#D�:�C	�4�
�:���=4�N$T�>;�;	O�����)0�>r�����+B�!�ETz�gS5����)/$P	��&��d�;.?�;�B�� �^�_˲anL��)R{�[,�+5��g�..
wSn}w5F����9�:���u�q�%��SV��Yw� �,b1P0���r%7�&�I��5F�uZ\W�����6u���3���4+�76��,�p��O�C�H�x�V��[�>0?sz�Ze8� S�l�jh�v�@"U�Xw�����S�Q����g{a=/�}���É��R���=Δ�/\�g>�`�s����Y �_���.���氂>L�ý�r|~O������d����Uo���]�+E`��E��@oյ��gJ�@��F��g��!�BWz��L��m:�6�~�I���
q�H�.]���y�ń��v���N�����y�� ���/L�0}`� qD%z��,�r|RG�\pĖ7���yN��L��˴J�T�ӝ���)�o^S_F�j6�����$�OƎ�B�~$��E����a2";��T˓�,�-��I�Gx�b���i��1U[�d@~*��Ŷ�wM��gU"�o
����T%�O���F$���	������y����'���e�|
^�߱@������k0/x#<�g�}�O;!����3���e�0r�I-"���/��Ί�3�>M�֌��>��r�,�;E���O�^� J��!�m�mï��Ὧi���䊹���W����RԽ�r���/�%��^�d���v���K4�w�n���Ga�wX��dH,Tt=u��O-_Uץ�����5v�l�.ߐ��X�u#{UF�Y��1t��'럯���:�T��ax6Y����!��Q~�`�	�1�٣>�m�Ŝ���j{;>�
Ψ(�;g�Q���t��D�^"n�2�V�}��1 ��Y��VU��a�yNJ��(ލ7��V���5`o�����_Ƚ��Ӻ Ü�rk�0f���Mp�ծ��U��2 ���jK�+?|HIo�21�G`� �5��}�Ŀ(J~1��I�m����V��j7g��rY�|2�M�s4E/����#�/���8&�4�h�|�xV	;0<�e��4t^H#����Ǥ�)zƫ�ٹ'Rˎ��o��!D�T�����_y��S��&^ܶ#д�%�꛻��7;^�`�V�z0Vy9^�6�uou�rj�]"�(�8�V�V؇�1��������}!�s2l$�,���ů�x���}%q%�zl���*�qg�>vr&�i��[��5���_|ഉ1��U��&��ZϠ��� :2U_?��� -���	N�{���ݯ>��?���'��~Ǫ��'���A����E+S�ޑ��#�+�)0{yJ�n��%z����8�����x@�p+��ƿ˹\����8p쎎6��^4�F'�w�cO9Į^�cr�%J����^�~��vz.{:��f��9�St�J
���#Le�G��H�6z=n1��o�`W��+o�g��"�<���F�[��;:?U�� �˒�|��SRxv�y�Ԭl\R�AJj���nN���(rPG`ަ4��p�ʤ0h0��px�6��§�`r�u�����mv�N=����O~�)r���e,����.a�����O�/���W����m�@��3K�W]-١»�$��ړ��$r�nm��B<��k���'f�إ&���jx`&�_�R	݅ ��٬`�p�C?��=T�=*��$��.Fk�"��#
tJso�?9�j�y~\��YX>mR�i(�ab�A��� �~�����C��9,\�t�)���>+bƺ�F0R��$���+q �����Ҡ�!
��6U��i���vI��Cv,L�RlU�EK���X�e�o_A�~�>6�ŏH �Ib(qTrI�ɶ�FX��IR�\�u�|�x�ͥɁj�1�-�a����h:��������,k��AP!TwUP�"]QP@Z��J��KG�zD� A:�C�	=@(�|��Ͻ�����������9s�甙9S҄�{�|e�A %v��=3'<�9U�ԒN|ќ�nM��XbہK�ڃ��,�ӑ
�w<7�6�׮�K�~��-��g�v�Ս]0fgVQ.��{U��yt.� � �w�v�h7u��R�9�?!�:M�=Q]k���ء��;��� �(�� LYP%k�|g=>J�ܳ�S�0�a��8>���p.��=�õ�#ůY����Z%6�F�Y#΂�Ne����<����u��S��L�nt����5�D}݂Șm��Ր��x�{a�r�ܿ�V�x�ᖅ/�v�J�]����h���bz{�Ҿ��E����
o/i��������H���k�;�}Иn�Z�oN�����8Y6��9u��=�W��c�ly�ӎ<ǀr���3~0:^{��Pm���g��=����Q^XF�.W�����~��ǈk�+�aG�8֒}hkMT��s�w_�MI��m�VaQ)z+x7�Oo��Pl��q�O��W��6�ї�)|V����a=�l�Pva
��L�-q�#��)�{R0\�@y�Yb�0x�u�E�/�i�#i�|�k�b��tJI%�RC�?w�^Xn8��|*������'�-�?�e�9<�fR$4�V����<������y �Q�%@�q�Y�'�k�d�W64[<����ɡM�eȺ|�r�E��V��W>%e���y�:yczcF4�����.j}������n�31}5�,�X�d#���
�!P���+o����ہt_:音=�]68E��ˌ()�������<Fw�^�8.o�5��:7ݙ������K���LuV�_@x�����{��M��aj��⮶��m�2_lG]�)
�(��	�ˆ�alR��#r8�:S��%)?:s Ko|�60�m�۟-��w$��b�#:K�M�MIzs���BӡBߵ���=p?�N��`����� ���8H��j������~$IX�n�\<[���}U)CX�'��e}4T�Ua$��@��I��mo�M?�W�Ś����Wjn6'������IԄ��FX���f2�vY��>z=-C�ֿ�hH�I���;���P�:� ���n��Y���ys���7cx���t�E?/H<	�P=_M$)bR�����HC_J#wZX���SPJ㨚�a�v�!\t�"C�ѩ`�t���3.S��+��!�}1ݻ�m������lA�g����O��*Y��Vj.��M�I���P��R�;�hv��a�f���qC@9[�3����?_�����)�O�B���2�-�b{��V:��P�g��a������� 	��"��7�F�ﵣ%���_��%-�</�s��X�әU����K �����8���A�J�Ջ%6j��T�R;�]���}�겂�<*��[��I��sk�U 2z��v�7G�q%H;��(	V��K:}zEtRoo��8y�;�Bi*�(I��g���w��/�]��~Bۖ�f�ҞD���G0=�&�[�.)u�"�.c� ^�����$�i��@j�M���)_KP0�gl\g���iEԶ���<��9q�w�R����'߶;��k�bt>T�y�|"Q��8�B��E]���9f�ze���4��V�)�#V�Ћa}b����(��.?|b����A�ɬ��ԑ�%r�
�(�lUGR/�E9��.ٚ��y��`LdfNE�`��>��RV�>�U�M�p��M�X<�j �Y�)���6���o�&�0#J��F�MS�eE��K����4.�g|"099y���%[I�RY1";u�'�}ݬOW��nʤ#��})6���,��V���>S�K.�k��Зn��􆧚q^��.sX�qFb��p��~L9R��3H����k|�m�<�N҇j�jSw�l��Y�:��-!�gn�����m��E��_hL�Q?Nv,�k�M�!���]��=JT�w�?~����~�Ѝ�dy��*_�����2��v��-t���Cw���V>��R�^�a(VD�4�Z��]H`@23�p=�v\I��
�._��JܸW���γ)�����i���b\cLL�P�m�����=9��X�
��E6v[me<)M@J�^��Q\�ѣ� ��~~���ZL��5�؂N�ϘN����-+<�b����l̢B�{�K�;)ʊ����|�ϗ�{{{ێr�!�h�u~t��1�.�9̖p�y�ISt�)y�Ҥ�ECc#2&��C�10��{�j�ڠ��_AW���rx�0~-PIF�L-ʊ���~ඨizL�J��O��߄y�e�~�|�ZDv��*�%�:n�Z=v�.�-Mb��!6=�ĥ��g�2��vٕ��v�����Z�U��T�E��^��gWl�{�J-�s�����"�Ss�,����ﰌ��mD��aiR{�����N�T���-$xת K��z�R�Я�_O�×	����XI��HF�y�=)Ob�
Q��UJy��<�*���G�N�K����Y����j7!�R����V��0�;v�x�R���T [�`���d.	���P�fj��]�c߭��?��,V���������,g�lҚ�(���˲
1�mé@)�'�:/tf��z��ݼ�������̃�qq+Þ���������(���j����{
R1s|m+��a� :�<f�Nuܮ����!�Df�"8���W���~'��a� 6�ˇ����~�+��B5�Y�u�nP��ľ���N���(����OjM�I�9G�@ny���&�`
)�j6N� bj���t�]|u�E�L~+M?�l�%'w�b�'@SRT̗� (�h����*���������;2 `����zj� * d�v�i11��:�u������'��6%%'�*�d��\X�Y)�S��V���~�\3���"���@0� ��mT�d)����;G��TTT�f{r�w(�>�<6���c�$�e-4�!��e�j�u����u�]�����Ri�-�����1---�E˿1��z!4�mj�>'��6� w�yH:|] B ��(����4��~'��;� %�u�
�	;�"�1򷳧�[�s
��iy{���B�ҕo�k-PY!O#��l �-H�2�ӵS�S@4q��an�KP%����2N� �̚��Ó!��7��Eށg]��3՜�Iq~υ�~ ��	X,�y�Ɨ���@����]v#�������_��� �}��J�j+z�}ez�ʂN�a/�$$�iX}�O�w����d�Ӣ�dM����r �Gc8��ٯ!��.�����_��	�Ċk<�Hŀ�7���5�%P��,�ɒ�~��nw�y,GQ�^f����ߎw1-mhԎ]�z��`@R*�Ĳ]�E�	8z�x�I�w��X�S���o�j�:�gg�n��o���
�6,�ˉ#�ހNr�~�E ����t�t�����U������\��"xSy���� ��q8������v7�����I�A
P�/��-���N�ϱƗ�rp�q ���#K� U�������m��{<d�o�h� ݪܴ�yW��~a�:d}> ��v��@p�5yZwY]��1�m44{�l��a���i�D
��ޞ����iu�҂���֌1�;��-d�
f��t��n�o�W��ٞ���)�)j��$��{ZZV����Q����Q�ee��s�v����ͽMH���אZ)0��s;�L�4��&�ᄄ7D��9�IK�����(Ah�7��HڏݎE8����}�^33775������	��V�����t�?���n��.J��`�1����� ��m(�ܞ������FUM(�{�!�x'KP�����k�#��~�T<��Ú6��F�d���~��	ĊW1*���Ħ���X(�.�HC)�E��c����\��8M��A5�w��FgO=��dTP��6m�2���/(n4]�����LI鴨	�U��&�]BA9��ʏ:^�A�O������/�Q�8b+�vnJ��K�2���������2�Sɡ��8�BP ��2�#0� /��h��j��>���SIzJe��՘fh����/���اW��z�"���N�+��?C�+�m��b�9 ED7�G�H\��(�6F��7�ܦ�����v�C�Pi��|�d s-��a�r�E�C�\��ֻO]�����/d���n<謥���*����K�$e����Z��%\���6AqǾq�G!t�!��yw�	�|�Wfd�S�<��9q+4�N���f�MFW�G�:�?�T�}k��u{�4�8'��� ����J�&
&�=ؕ`��9yy���S�n@A����G�Sz���8G�Yo�ԫf�h��@��h�kV=��_��UH�'��r�H��I�s<k�lKb�:��	��(V��CG��b� ������k5X��J9�?����JA� �*~@U��0.{�0{4�}�h2)Z+��t�ڻ�C��淎�yQ�2���p5p#��h�����ڞ�.�Az��
�#$��j�`ٮ�DC�+�޲�v9%�<�H��S���Cϡ��8-��Ժ�U2�nh���e��
+�P�9 �@�߃Hw ��{�@�����d�׾s gM��R @&� �A�nfvncc���!�)�]�����B����xf�Ũ)T#nGq��)�:zX�[Q��η��s���x^FFF� <�B�y�j�uc��^�����`�ߏ��u�W�X�S#E}��4G�>4feʧ]'=�����fv��q���2 �����r:�
�������@��2#�p9�W��C��@�wx�⏸ot�B9�ͣ��}�[�P����d�V?($1�Z��ʖR����p�ii��ܦ�2�g:��`�F,�ɪr�O�Rq��7�Z����9;(*� �5�-]ޑP��Pf��>"Pu�-4""BY [������8�TB���Y4��|h�֮���ܮ	��Šѭ�:z�ijiힽ���bfީ�mM���+�r��kK��T��A�y����J��zKo�R}�^^.��]�NS���O������F��*���f(�� ,��9f׿%<� �VXq��2.�M��^%F�-F�k��q� ܍K�t|���S���q=#ʉ5e����h�*����p�w�d[�-B�$	<���w�j��:�m_]cȟ�4uɱM1vhҘ:Ek������L5N��8�CqL뾄�ⓢ--�X%�`׻/ْ.���,�����S���`�ssj5���T3h����@_d��r1��'���/Z���Ũ�S��ܵ>��r������D3��]ŭd�����rp�n�S����"bg�h�U8ݮ�͒` �*/kl7 �_���7ٿ8N�����H|��:��Y��<p�E�h��Q�}���<�)O)����f���/��W�rpqz��芦|�f ��M�_�e#�s���0=p9�ec�4�<��H��}	C��nv�ck�@��;��8��- ����Ui: 3�|�hi5cLķuw�̓G�@xe��9 N3�H�.]���/���Y�?�H� ��p��Z�IEx�Z�0-?~��������a���i��1�?�D��WK�b�+7
[]{�f`N�����r2e��!�/��P�w�Ö'v8�5}[>tmt�V�i�ss(�x�N�|u���/�"5����#�u�N%��;���Ϝ����`iD;?�t�d������Rk{&U"����{���TP�k��[<����^������D����lJ����'Ų�Ϋ$�y
�U|�H�M���.V_�,B��.[H�s��X�l����g�6�����q�'��`aM���?U��ۊk߮<U7^ih�'�Ғ�0�p��_=R�kz���x�"��Qtn���ץ� r!̟M�[ګ�2�Cc����"z��������W�/ˌ"4o�ꗾ��]��&���k6겭�}�@��,�@��Sd�4��8�����m��zM�Ym2u����9����>��������Wer�Z�I�T��/�V�f��7i�C�-qdKf(m�j��0wf>���-�sಜQ)]w�.�Ħ����t{5�k_����Z��R��;�8�j{{Q�W}���a���ո����&{ٛ�`u>j��R��$����FX�����B�\9!O�?GW�V�g$�Ό%�oW�7�M����V&�_���P��A�窹�KWsf���K֤�p{�-�$
I��7����Pd��_�g^�J�\c���|ܒ��#�	'���+�B�0�}z\�*(D�m���nSg*�KǿMn�h��4t�����Z��yL>U����+�1�zx��uS�ZQ�!���Bq25�@!��v�>Fjj�� �5|L��mT���J�[O�' diҤxQN��\<�̙��E�G��q��������V�Ul���/y-�3���(Mk�Lq�M�G��yjx�s4�D�J���P^���@&�ңfF�މ~�s�����sJ�ǂ�mmtL��#�褠K�H���W�=����e�]�&$W_�����R&�ۑ���%�q�N(@z;&�`�3�[��n�3>��I���An�����VBԭ���S�#���j���}y�2���Ѭ}R�@;-_L��/���K�סg���{R&�?����DFW�p�����-r�E�5N7��'����\F�	���~cܒ妮�H:��k��s?�}�+1�<Y`��*�[��^�?0�X~i۲���)��>�]��������7�%h��r@��d����jbέΥ+G��[�o�_ q]���Cȁ�������!�QZ�pi�������Դe�Կ;u�+3�Wዑ}��ܥ�B�p����fmog��d��|���v���c!W�
��[��ǣ�"�Cy��ff�)������h����J�ϥ�#�[R)1)lpq8Gu)s-9v4 Y_��l�xj>p�Le�1���Ӽ(���EֆS�&��Xڵ�B(��kے<�e�cM�cw�X=<�5�S첤��Ի�bn�����O���l�)\���0ԨR�LگC���"�/) O�p_-���|�.aHnً]4�a�{�7x�D	�xb�܌���� �)��R��d�I궃R�B	��>PF��Z_^|3���������'*W�8e�h2�@����F�����te��/�{�}Ie�4eU�v��mll,3.��]fI֔�R�b\>ݭ��$x%ELJ��[-læ��+�HI�-���34�f����=S��Q5�QS��twN�sc���~tl�������7�N��4����N�u4���z������T�����^����;ȁM�`wc�k�m-�mx�&1�����Q����35����2���b���JA�� Cp[[*�T;|��4py;j_l�o}��b��B���e'�������)ug(y�l|o�[uOᩀ�[c,�rB�kn�/�O��i����%�G%j1�}������������L�%]�!9WB����5?_W͛���}ɺ���R2�;7����P�©�h��R��9�b����^ܤS��@�A��8�fi<,]����XNv�Y𝿐O)������P�	nA��LW��[�uF��ud��W����\p�"��� �G.'\�,&)3�ť�U��	O�隭�W3W|��!��q'�SiZj�0�d.��(Q@�J=X�+��lP���5�
\�u�#��ta�Tfwi(/��R����v�K8�b`�9�@�_��Y��z����E��������7�ٝ9Z=�m�bśT��#k�7��3V��XY}Y*�j,e�Rڏ�plC�����]����>���z���Pk�x��t::��b�ht�\_Q]	!���d��{Q^�����[O|^D��`����ތ��\<L�/��c�L�Zx���T5K��+#����Yg5�ð�F�&��=��.��%����וڛDb��]���9��6A!k[�KF�������aכc��[�q}��	=j��E"��aN˼+����y�D^��+J:��D"
��F6f�A�1�2��E�Ǻ%0`���FT�/��P&�]g�F-F
���fL+����}�����J���)��6B��ySݞ��,���*�0D�E�uԈ�r293���m)R���̠�3���>E}�H�N4ǘZY	w�����30C?����%�b��������i`���	;M~s�ŭ�g�Z�ϟ��4��Ͻ�_tp.ɿ���'���6vI�n��<�+��v�ߝ`��;�+�A�l�纇?�f�N	�K1+���;���q�^cZB�= ��k��Qʂ5*F�!km6>�t�\�Zy�6	���`��۾�����繐R��W&A��VT��2��w��c��b�2�m����ks#��wV��x�M��`�'Rja8e�@�W�����Ny�-xY����y8�,!�L��uj�8,'��uL��B>�^�Ⱥ�!�/�d��?����Ny�0,�5P���@��`P�������> }�=iǌ�uIS$RP�~Q�n�G��s$'�n<pxOE��R�$7�h�8��4Z5CV�Sjҍ����.���i��^�3�~�k�6k����Kͷ�y޸��@2WV�|��9�g���$
�s+��_%e��o͚�Te�
_����
�j_�Mzgm�>#"PwCn�=�|r���d���x�8�䳸K�A�=�oXVȊTn.R�(��~�lՙUd�/-��mYl:&Rlҙ�(=�*4H�#Q<�w��J�փVj�7�EQz��%$u=���]���Tn�U��Ў��������Z0���b��[[qLW��b���vB�<0�^��tUx��GX��������4T�@fm�%�)����ׯ7�z]����^}4Z`7�D�q"ı�;���@�q�E�2�p~\?cz3Y���w &��0vJ����EZ�Jy2?����6�}��K�F����Z]K����ʛ��638#�l��/ij7�c�כ�(��
'��V��q��G��t�m�̨���?����b��$Y��9>(�,k�����}>J�e01�/��w�V��3�֧Wߧ���-��;uɖd(�2�I!�N
{;Vq��%i::_#�⸲x�{���~�z]@
^�B��l���� VOB�nm�����l�ş�)�u�W>KG�
��)䭪����n-⤭>���
�B�~�
��#�B��E��A�������cXK����S��Myt�:I���*��|;�Ⱦ�~�P��5o�=3�_�<14���X�j�N�n�fӐ�8[ t�L���_r�3��b\
c�Vb-Z	�1'Q��J�x�d닕�־ZR)��C�u:H��/8 ��2x�Q�5w[�t3O;j���Lc۪�C�3�k��VW�+��C��X���ӂ�����G��F�͊n�O �[�q5��w㽉�%,D�س;�0�"D���S���ovt?�3��şj�e\��_�D�i�Z�#��e�����~��bR�k);�������{ G�!"ͥ��ovQ
h������Y6�	I�{�T��w"(�}ޑ�
I�b��a�[[`��@�����8�|�z�l���>A��XoԌd6'$��R��gx�bNp���[�q�Nh��<��A#��3�,��=��u�^t�yFY��40�S��Sq�렌��E&>�Ĥoԍjiűa"��'���Y�#�^^���uY����0������6�l�%or���y<�!�ln�n�,�gW+�m�n&Y~N�R�b*ێ��|�ہ+�<U��N;��)X!i!���_��Y� �$��&���.J~��n�+���]�ܿ1�cNx9+�D	܉�T���O�8������_��c��b�=����s�9��G1�����֣��JO�����3Z�P}'��Z�S}��cr��䁉�/l�o����t����Α+�mY�R����٧�����,��[�SG��+�R��[y�� l^��.uvypm]�x�A����{�?:���l"@~gI~ga����n�o�p=���*m˸��L*�������B�Y	\A<����8��"��^���\�0�_�8������I<�n��|'�I~k�L?�VQtron�1bK?GzX+��r��ÇP���^�!�ԝg��[��7���C��Ҷh%�ytE��te��qU��v]bRX�d��kv.���y�ܲ�s��cW�E?�</��!����ӊ�;�4G����u��nѼ��͆2��E�5y�N��ݪ��T��]���U5�����<9�CO��I�SYd8��^1��G;b<��zfk�fk��7���fY����F��g��r�zK��愓���+��'�.��,���,����Id����uu������D�(�B*���~FcF5[�h�-aΦHіԔx)���(NS��;�q�D �CS�aY�����;�esVO��L�`a��,�-ϝ;��2�a���a��i�ˆ�Mdӎ1���T��TL�O������9�9<��S�ɒ�降��q(��7������VZ�b��.�����y�= ��-�����bG��Q�6J��F�����L�=���R������X]���#1
5�z36܍���U�ny0�,��Ef� �����P8e6����,z���!A�+j�o>�e��C����B�̚�g��|�@m���^��������xL5ή��A2KN%�G�����d��EE����`�6�Ʈ��ў����z���E��%"�����:	̿�aeBE���E��X��S�b��:����EǱx?z9��P�O�E>�ϩBNƺy(mKN�l�#у����><�w
P�fU����,��[��77��ѯ�${u��)zM�F���Λ�e����U��G֞��=y��'qm�G��j�1|��ݠJ)ʃw��=�[AW���A��TU夂���[�.�eơ�}�zJ9�+mQN�Y�U�ם.e��O&G��ŭ�Q�4Yxܩ���L�V�K1)������I�����,��'8VF/2�!I�z�Y�����;L��`�L)b�D�w!�pH!'?u��'w�ɕ��-ɯ�yI���q�b����W�C�~��6�I���e5��z1��֕gq>���Ք�:�d$�7S��}s��2b��u�F�p=J���md{�LA �`7ZI�<(��� �H(z�E��j�����[dWQ�ѣ��$`�0NS)@��Z��`�ԕ�u{�6|.�ol�LI��JM"��-]�_�m�'����	���n[d `@8-�*����-���`ƶ6�pf��"`0�������?�7��є�sQ!y�+��KeOi�lr4��cX�3#���Kfs�j�tė��ڃ���z���&pO�r%�}�.���󐎽o"��<<P!qJx���[z�RS�^�U.f�'</f�oq�56Gu���\�R�nvN���_�7��a�q�������\��b�ݳ��L^9���ᩇ��~x���!�W�ttI\��?�z��6��/tO��TM�;���G�6�Y�ҳ�9
��D��O�����@��_	39�����%���%��7	V�?�_ �?��$����T�'�bމ@���%��7V��̂��(��������@��������+t}�IHHD��:�}�������:��0���:dc� ^����A[�g{C�+�n�T�����5�L8��r^m��*��.�DcV�OL/�K?'�z�l�?�3�yl�������5�����ݠ}����t����x��H�[+�*B�bT��ߑ�_t��N
	B\Sh��g)"�)����Z>Wd�4f���>�m�j����318zd'B�%��ܞ���W��-�vE�^�m����)���ĵ�L,�Z�30�W���U����[7����������P����е?E�Q�\q�_�ɑ#�j4�W 3��@����ϴ����9�Uֆc9e� ��;ۄO��c��v}�����Q���o���,kY�M>	?��`%;��y
P?��gg��x���(���7gnK7�t!�� l��J�=˔�VM׉�6�^�M�ߤcd�7���=�7����|GHdJf�p4)p���]�* �y'�V�'i������URQǎ+�U(�Wg���A[������9�}��y�v�c��g/��!����o>�m��㧍�$�k�kM�'n�m+l`&�E�=�e���o�1a�hi�
;��,��K�m�߷��+�ݤ-�P�_Q�\���W�AX�.������H46�x �{G�6�#����l��\��kS�~�[�� �m�q4�%��+��$����,ƙ�[�+�WW�=���g�-�r��A{�W�W��_ �24��ĹW:�����}�&赯�݊o�f��u�{����0��j�l���c�V�m�v�����ـ�7�e��B{{{�~����#(�l�o9x����ݰ����{FK����j_�҉�f�s���j�V!�J�wre��reӗt��f��3t���D|L���4����/�
��V���mJp GPh�� �y�����b���G�����cM�i�=� ,�`υ�F�hj"�B��?�V�ޮ�H��Č����Ə�)q�.��p�.�S?a~m_�S��\2���lZ".�/��=~�͗����9!�n��8œ��u��1ѯ��M,.�G���l�Udm�?��{�����oj���Ɔ�0aV��]aV�V��g�)�s#/1t��DG�yQ���`���F���Ƃ�y�� �֯�+�W�j��r>���@D�R�2���c�j�{�x��V��/�4T�bu��6l�JT�8��Bx�D<�F����1237?�^	���;�>��z`>�j�	�δY�4����5�m!Ci1��F�yЇ��V{�����6����p"�c/e}I����n�G��bݏ�V���z[ܯ�'�9l��7G��:r@�6�|���̇���\�&.�k�Q!_���rsm���؞VFdwyQ�lA'�qK��*�cam4�p2a����G��6���'M�ϙ���?:D�*n��g���ŗ��Ro��X_^
����xnO��Z�-"S��#��׬�r�zT���X�d�$�x�}�����KoS�,dm�����D�x��t�┬����D���1�7YK��GP�V ;�����vu�8v���$W�4b�� ���D�|�ul ��JN��4�͝�%��Vs��p�n���mZ��7I��ˀ��.�&̺��W���m��H�X���J\c9�0vH�MM���r����\���1ă��&�ܢ���ty,T}����ܥy�CWt�M�l{{�z0�zp¤!��u��CĤ�X>��b�`n<=�AB�ki�5}6�=u~�V�7�"�t�m�p����[���=e����&og�V��/�p�ז�3b��(��X�E�e�6�Jǔh��m|.hXr:U�HPml^�"n�B��I����X�`��N&6���,��_�޴�A����a�4r�.4�/���>��%�����L�|��5#ٺԶ��oG�d�EM��U{��������=&�?�y����/C1�ĿԶl�X��FY-�?��ŞjD���J.�=��g!��i4p�q�%堪�\�k�]b�#C�_��t鷓�>���*q'{����%#��^�j�p�ޞH	<z�/�8.����l9�'_�Q5��Q2l~ظ�ͰMS�Q����u�������F��C�6�������܇U� a=��O��͖Pf=fդY�>}?+C|�p��X��Y|�x����7bw�ׯw��K�.1���'�vUt�I��bTcUA���(�Bv�,��3Y]b���>Ԍ�x��Q���v]�a_}�q�p����U{��q|�ك��ǸMu.we�/�浜72̵��2k�'�&,y���v4��Z7De*�����b㔸�Ƹ%;lBq�P��ٵ�N#�O1K]/��vA<�)`<���G�L�8g
`oQ�:�?�p~�Qcx������Rx��M�cڪ��~��u2�y�O�|؝;� ���wF�u��<]�������s�7V2���a`e��U LL,6۸#��S�SSSV}��+�Y@���{p����ߛ
"u
��R����_��qȼ�^y3Qh��
�HNE'�w�þa��x7�R�B+%�bu1)��O8������b6��۞[�0��z)u�bOO����gb��HM�o�;����U4^%���8l0ף�g?��x�:��1K-�|{r�e)	�+op=n,	�yV�(�*�֍��Y�r���sz��7��Y��A�57����>�o�D�aм������֙Z^�%l�Ͻ!����t@J/�5s�R��݉]Qy�f!�j��)����G��楀�P�v��AT�c����]F�����*K�V[ .*�դ���'�k��b�~Rғ�Vpb�ˇ��kMV��4���ҿ`��WM��W���Ɵg�k*�]�=��43S�t��!�<f"�K�ؿB�V�7�X����o��6��Z������=D|�:d�%�_ߥ�Bm<c_p����ۚw܁@��3�@��~�ǟ�5��.I���$ޤ�D��R{����r	zx��J�z~���y�nLtKWjZ�Iu�2�G엣��,�E�1@:W�2�e�B�� �TZ���p}�t���I��;gk.��Z'�w��\tqG6�n>4������Y قș������#�1�~|:O�i: �U�c�A�!\���M���.sO��f�}q�&*v�� ���/�5Im��Ffl}�ٚ�_To��ӼR���'������\J�Y76��~�<��m}XʥC{5  ����mԤ�+����]�]�Ƶh�H2W���Pf&�I�g'a���"������-n���M�R��`� {����8�����Y@�Q�O�w.��x�$����7��ЉcK�S���	"�n�_g9C�F,���Aπ��G���0�'K�V���sA]���Pg!���4NG�>5q�L]��H��}�w+��>.Ԭ����xB���^�BW�U� J�U���h �ۆ~GI���8Z��P8�m�ץ�)E��G�ڞ5M�א���ęC�K/t_����Ԡ[��Nj�*�w[�aI^~�@��e�h�=�NMݲ�=�b�JϽ L�Q�3]�$d ����E�v���"��#���R׫�7�Dj� E"�������u)��Bw���Љ9ð1!�;�?��4to�a�����X��	H��]�փ>�µ�50�"�}��E.]9D�&��1Us��n�jІ�D�Xm��7��بǷ��[��7)M���D�Yl�.J?�a�q�ٯ�]H�����J�SV|������	sUe�(w�&N�^��j��1�g����ɪ|�wƛW�7g���i��1>�]��C���O:ޣ�R��*��P;�=&m�rn���0���w�p��#Zi`��.�ׂ�W��S�*�6���u��y2����ET����Ε�5DU�k�.�>��NdAI���wΉ���Q|�`�z������V>��1������M�Xlg�.��F���5#�X�N�H���ȓ��3�d�#�4�16�t�����n��U�����!��S˯Z��P���n
��(�+�߉��f�:�f5�\I���>d�*�Ib���Nׄ�����SY�TA~����0����̢f�l��NH�ӧ���v��H�q���TZ�w(�?�E�o�O,��tXo�ay"��aL"�?���9���!LO.Ht��Y&�|����M}W��p��T>�m{-e��ǥW�Dͯ����:镅C�����x0?���jML&J.7���cU����%���3�i���$_{�M3�M.���ۋ�|q��� MQS���M��x�k1������"ቡ�5~�G@���?8�JCB���6����%�.��A<��$Kh�^���y�ܼ�/��{���~���Cr6���v�w#�q����^瓜:K���]Ľ��	�����qM�sE<�u�?�j�Y�h��E�̷�n��%5�p�YnE^[n��3�����ƺC���O�!��-N������譡��a�f�"w��L�ݥ��,f���a�.����i"�-����l�������EK�ʃH��;u����N>}�F�B� ���jHX~���=y>�n>V���{ay���l,bMϢ�_���7dt��x��26ͧ^0pS 6��5�w:�g�c�(��kn��6)�x���3FFN�F濧����~�����"+�� ��]������e$�k���?��&�1����5Ɵ�:�7�*2����p_��QS���/h����Q��>U�b)�6ݶi�:�4��h��S�Rҕ`����бe���R�	�c6ӏ�z�o��gy���%��R^�+�А���♅�]��Į�.:3*l�H�ם���4��·�|>T���T�+QL]F���q<_}8EV;�]�b+0>ouqq/d+$6~�, �)�`I�@^��޳|�*l��v��d�`_��@\�sl�����WjeR�.���{I�(�%��V��N�BvB�̜c���C�v6���W�y8�C�?���#4����QO���2s)����k>c��Nԣ�%R��;���s���|o�֣��Ӆ�|5���gG!�������^%��*l�S^dɟIg�u���O�G՛#tN�.z��M��8���5��i����ό���y�ȥ�U��,>̀P�7�Ɵ$�[��n�
�0�*OM�5��r��ta���7�rZ��@W� ��Kw�z�DU�g�&�'���v5�Kd�E&= �! �dk��+]a��⏲�W�녇�t4�~���+�3��j�Vr��9�LC���Q�	)t��L����(K��T�w��/�Ԇl:͍sfҹe��E�WK{�BB7����*-���e&��'MԱO�ؚ��x�B��鉲��"�K�k������MK.=��p1���y�=����PH|hr�b,^��Ϲ�w��l�b�f6�<z�Oʽ��қB��$�Df�7�p/�|��s�;U�1���7h^��V4��?K㈿�������N�D�{��)�����_�5���o-_#O��SÕD�c�~hg�䢸�O���J��>��`���|z�� ,G6�iɵ����pa!,���P�LOJU6�������j��!�����&�,Dw�`�N�YE��W���w	�d���'j7oa���0A.�coKl�����b��[^qtc�k�@��LM��'�o���P��	�;���Gl:`����(I�e@)(O�]iB �q�W�>���K%�*�6t�~]��k�ub� ��;�����N|:�침��{�oU����'<q�$�T>�����ys��N�R
!}4��-t���Ѵ�
h�?�e6g��Z���ӫ�g1[���.B�B1��3|UFf#Dڋ�by<�K��B�?�W���3����d�M�����3a�	~�o�!w xh;�na��Ĵ��A�Q���)%�#W�`&Uǿn&�D��������MvN�R�U���G���Ն{��9!!K3�Wϟ��8�~̲{B^`}���j�k�d��>��R��?���y��Y%>Xq���pGy�j��I'S��Cg�*��D�k��=ZP7���L��\�^m��p��UH�%>D����$�������<~���#t,��U������M�	�$�B%�7L�p�5�����J_=pz�� 0����/��iĊ�W�v^R���,�nt+�A�Y����-�%��g���-�x��vt4z����[�~�����Z٘���2 E�*ݴ���o����L3�M�*J�և�ɠ��R�8�9Z���� ����Ak�����P_{Io�^	>�v�p'X�����������]n���m�L]�̤Ȭ�!�(SfJ����1��2���)���2Oq8���1��]�v?���=���Z��z=_�����k�j:\Tأ^/v����uE����R� }G^+il��>ɀ-,��su�nl���R�ŏO;+�[��[ ��D4�������s�8z{-8賡a�/�>���~
x��$?�7
NF�rg�m�B6�=�iz���Ʃ�����眵�KtZ
���:E����O5=�dm'(p]*�H���B����ss�V��E�9��>H�A�H_x���I�s�}�m�Sfqc6��/o����C�p���J�u�����=���/8[�_��-���P`>�iKp���ε"�y���`6!���e|J{z�ʂ��p�ιy~a /!]���7�[�c"e�/6���(���?����Ǩļ$��-��+2DL�u3P�
ޡ�/Q���z@Cu�V�iH��8�P�{X$Tۮ��?uj��^ps��[WDO^*��nN����%��C�gdt�g"��/��xC��E��%��B��S����ŵ�z$C�b����0eu�9��\t<����5�=g2���+�5�/��3��e�9['a5�G9���7�뀩��.ǧ �O��]2�هac���8h<��8��腂-{���.�=6%r�oo*��"�2;�C���E�J���Yl��6
K&�;`�=���f�4�9kE�=��}��>�rO���}�<���	�R�{AD��e%�H\fy"��ۄw�f�i
�E�梔�tv=���~����}�zd�^�i��}<d�5��kg��Q��j�=�{�P���0�6�1��lW� ����BH�3�����f�Z�>���s�%��\	�Ǖ�LOd��ٞ���p�{J|ieI���5p��Ԋג�UU"�:F#�n��쑛��[?��'� X�**�p�O잷m�z�lA�k5�D/
T�/J$�+(�P�J��Zy��'_v�fХg
�cQp�^챙"�^{]��4Z{IDi�t�{�^����uD�v;����K he��B��k�(3��O���}�Xk�[�wZ0�(���[N���t��9����4?WT�x�7��E3��)�tW�_^�$-~/�����U@;B8�����ʵيhx܊����,�kU�������mω��, g~��lf��"Ҹw ���,l�QT
�$z�~��r�.$P^ ����߼��U�C��\��ֿe�0ف��?��d:���&�m�`2hǯ`*�⬿oL�!ꣲ�u����R�ZC�ݲU�v��Ր���@�\b8c�
��F�}�� �2�q"� `gO���$�y�#��y�=����q����:�8g�`�t�.t��B
Ȋ��S��4}�F1���6����HK�ٽ(W��W��c�)����n\�iȗq۬��ת���.�x��g(7���?./=o���b��)�y���R�bL�	�ѡn�۟���kfC�~�'��S#��p+Ng��Õ}���z�I9��?��^��U�2�m���1P���=Z�a�l�	�:��>�Qt_�G����P_��[�Z:��ON���qe��G�p�^ n���\�9R�]Gmi�V�ȯ.+�ߡ�������V��
@ș�w~񫋂�5�����{�G3���c���{���V��/WdB���wVQ����"�h ǭ[Ğ�zY���(�u8S">E(n[fɷ���Gr���B���aZ)H�N+6r�R:"�e�F� �W	u�Q����S�6�V_H�?j�|��{V-(N����(��:�|�\w0��Z}]ۺ�{����#�a��ur���z�	��W��4�7�)�4��B� \j�Wj��7^������J�θ�<�7���x���p���V�>���.?��u�
G�2놧��!��;��C���+�ƕt�3ٝ]���
ؒMk�3�_�M����)pq���Z��E�U�{	ɑ����Ķ)����dm5��h�-Lz_L��b�(���/N+��+f؂V<J����t��u��@/9j�DWg�����%&��D4�w���V����t�1�l����A�ج]���S� C��)���(�bUT0:�?�
@[��+�8���e��3uG��u�6t=�_���N@��^?V2�PI/!�v��0hX���솘��<��>gJ$��h�����eFھ�%!�G�&��R��/嬝�C��O��4/|G#m����i�&�f�D��^o�=�A��ske�c9�Iolǣx���{jq�=���9o��\�����'�,l|%��� �[�@��$y�������L��E[c�L	�;W{Z1䱃H���3DM��i4��1(�G�bhf��
��x��x�� \'s� ���G��Y�D�H5����G���Wq��#���"�#їP_�d����7� �d��X��:�~t���p���E\�ФsxFF}th�$8���7��7�e��:�Yw�� ������f`�&	�˷;`o2OF��X��� -��8�}�$)���O*�H@��HM�Ϙ�J��Ģ�w ��:[f��E�����^�HU�z��0����9B1�S�T�#LLv�{�U�lRT�#$�(7}�u+���C��N�Խ��B�b0]��JC~�M�C޺��t���Ǫ�[�#㵊��ď�3�(����S�ſ��eS`F�hҹ"����e�Ѽp������(
���	W�*1��v�`�gR�X�������?��� z���gT���L?֘��T��m��B۞��v���9G��]읠�5dzFd���`�������͚@[QB�g������A���M�a�#��"!�P@���ܜI��dQ\x�F��.�f�dC�J��P����]��
�m�����������;�.���iq�yQf���15@5[c�rqT�hх˙��J��c���t]����M��w��>���\�-� ����~��n���`���E\�*S *^�6��-���:u�L'X$)�ג����}�K�q�;/���/�
��"<�yzgBbz{�=S�E��itz�[���V1�r�U�2�7�1��:�΋`�P��b9;��[��Q�<�Z^��9M�vu\]�:���W2�]5U�i����t�������	�؃P���)<��`ke�m yF�K�s �_�멿�\�c�t�n����)��vE��??��`�ǵ���ygi<^M����;�~7��)�%���9&��MpI��,ՃH0���gw�:����'��ǟ��S5,���sTM'�61�-D���q��Rcop��kQ�
FwzT0=!�v:'y{$����Դ��w�=��V��ơE�����^����_��U�c�*e�m	-ά��D����m�TI�cO�����n�	ܿ|�ǂ�b��q��s���l�ڴ�Z��q_��EH�.O&����v���w�4��7Z
f��D�l�#/���}N�ٮ�U�:����=9���-H� ��V&��_L�l74�����d;� ן�+\�5�9�]�¢��\�b��F�\�-U�1w�	��aDlʚ[��Ƿ|d*��i�����V�8��\'���y39~�@#�'fz�a��@� �aH��J��M���7��M2{���-\��70�����=������,�3I��nR7�I,�,zn|
�Pe�����/��:��ͧ{�VzI[Qwn�jG�Ʌ ����J]�"]��T���I��7�+<��(1D��\�D+�NG4�L�%^�o0U:�����P�������E���3�otB���@�9� �B(��жD?U��õ��`�gD��o#�d����0v\21����s�d3�����X+�QI;k8Bޜ&����ǳ����e��y�����Ƙ���vXl����E9���6�����va��7�=��2�Bv��Tߺ���/k��\(�����%�6)�u&���{{cv޿�P��x�o�_�(I��r��??Pz�[Nse��a���^��7��3|N�<� �g���!Iey�j��w�B�'Bb����ph��+�Nx@2�����,T����f`�����â�\��|8��JKi��n5qä���i���UT�CEa��4�]"lP��K��V��&S���r�����AY���7��I���	�1��)�|
K�����3�an�>��2��h�3���#�'!^��U���ij(��E��;�Laz�"ӳ��BQ�]���A�)5�L�s��T�Ls1	����m�%˘�N#����g����4~���(+8_t�V�\:uL�|2>�=�3��	ix��K���qm̔آK��;8)r��3�ͽ�M�~�\�'xF�̤E��A�+7�L��kU��sʠ�V�ߎ���{ul_,�]q 7�\�E�hZ�T^f߮���ʩ&��E�^�,�ߴ���S�f�ה�������>$�n���qgS�l�-��g����N|�}Șk߶�V�DsE�����*Ԫ���?2/�;��K��U��\jy��'U3��/o�o������:�&��R�\�RK���Mö�k�8�v����H�� ?T(rf����wiwU���[�TF�И&�9U����	*�����d�Qg�DXP���h�����DC͚���:te����3�ߓ���:v���󫮮�l�ט���:ԕ��u���8-�qӦ��@�4].��f|NĦ�*s8��Iz����:F��xDԔ�6���hb�$��5�9�P��b<e.�@��E�[uf4�*0
���s���i�(d|�w)�M�dwM2���W@)���?�#�e�ܭ��[�)6j���ޑ��a�rc��O�[uf������K�D޲ �e�}�ũwʫY�����!w.��teb�_mX�� Mb���W4�5�9"��֝gl]iۑ� ���A�)�^>G��Z��T6`� �zz���k��xv���Y�(�I<��d�fd�P6P�Qk�2/�y7%����:�:]��Q���ȹ��R_Q>�z�Ӱ�N�~�wJ��s�ߍwDT�6h[\���I��ҹɎ�r���m�ŖE���v���;�T)�X]S�]���vc����#6Jr��dȼ`u���G�j�gq�	�s�|�C���.ՓB��NS�EYt�IQ��!���K����q�(��W�s���I����7�j�7����������t���	�^���7��Ê��}�pG���)�X,w�$�����r�^Lt�pd��\�����ƙ��9$����̩�+�U����j�UD�x�0d��XU��g8Ը�0�����[ID�PL;�_G�#E��sS�bь�A����X����Sv� ]�����v~����wV1ErHk^���n����đyCMowJ7ݠdr�I���Y��§��Fwg�W$�jU�=��dJ��{C�4���}NQ�'�����i��ɚ�}�7����A�3K3p���e�L��c�_��z�0��UDG�ot�R�+q�f��$�~�T�����^0֒��g�A����rs�m��߱��w�����3{�
,n����P�"��L�l����>��t
qW���w�,Q��K"���Esi�h0�	EKE��p���韓��z
T��7��g�ly&Ip0v�_��Z�Q�jqn�7/± �9;����܆�O�[��K��&RHA%�wy�1���l�}�O0k_��'΋-���uE(��T����H3h�|�1#���ct�|˹N=&xփ\R4(�=��1�1@�())�P�gn���մY��0²��cPl�Fz�Q�v��}�fp���3�jȷ�+���7��l��f:N>ʭ�-#�HK٨[����?��a �WO�U�^���-~��w4	,[��&�>� .�P
㩅���L�����嶫T�T0��*K e}V[���"a�5;KjP��d FW���㒊����ʊ�Y�}� {�㻼$��(n�lw���%��C��c�ؠ\��p�h[^I욹HA�����R@�G���3��Ӏ�$�����okdP_x������ۊ�	�uF����ϩH��X�(���3.��sUvQvxq5K ?1Q�+�{I*����Gs���ec1��74���.�������^�MB��A��1�G���RI���ސ�َ݂�J$a�ݸ}C��~iT�͙��u_�Aش�hʆ��>XpndxRu2}��0�Z:��y�����L���Bx����z��*������#Ώ�F� fB��N����_����R�S[��J�DP�+�C�|c�!}wBz�']�zPV~_���K�:�AeX����*��}���?�+OIQ��=p*��
���Ƃ�f�B;P�k�����ϝ�����Ef�~e!��e���7
�������:���I���=*?5��ͻ��t'�#4���B
�go�l�>/*	G;���,y*�����ցf�7�[�� ��j=J�%V�b�=��ѧ�J�v3��1�7܀37H�Y���ɱ|���**8%%e���|9�[3PBd�spi�N������p�|@^cb���4&�36����Ow��磑V�&��4_T�L-���w��|u��&��~�h��^���UZz@�~'\,Ze�7/�^: �"!w���ja��ĲE��'^�����Ra�h��d�qʫ�1=�S��B*;9w&>����-�7�x������=xAv�l�3�_�א��:ǻ��X[��P�%LYǃ������r��Ie�������=��VlA��2���K����Q�M7����0�DWg��<��Qc��S�!�Y�߲��I�Y2���h+g�6�����E"���}�|Co]���"\l���l�5�����*�8A��gM�1����2G���_M�lp/�_�F��`�;�uU���~3�V%?��� ��dJ��6���c�N��n�ڜǣP�>��_��CD�n��-e^�tʹɠ�h���dĝ��גܖ>�#W��6����M�����FQ���_�ꮕ�M
�?|���� ����T�u��=s���|`�چ��V��v�������3�p2��W���V�$�Uy�E{�����l:�<��*Ɛ���(�A.~��WB��A�5j}ghY�~�1.���+�T_L��Z�l�O��خ�<��|�*BW݉�ο6e�8+-	R9pXy=�0��:������b�.[�OJ�脤zc��6����G���qB]�UNf�o��M���Ԑ�;6M������y!����$Ѝ�`�)%��5�a�?�:t���1�ѣ�I�q�#3�?�H�j�Ϫ����j�9���������ysq�5����aD\$��#��ɕh�V�.t�'�Y~�;R���S����c��T�r�P��{]s��������٧>"�?��|��v�ˡU+���n�Cԕ''���8ɁS�3A '�����d�c�P�A�s*���sm4U�V��K#��N������%w��:)L0F�oа4���F�Z��
P���L�U�M��s��ѓ#�O(�g26�6]&N0��I��5���?�!��6'?�nQ-�:,D���+��L_�X��VS��_���C�5E �؅B
��6�a�	�M7�McY7ak�Y�P���X�mˉ��K���%2vë��Нxi�0ߠ�|*_��(W�b�nm֦T�)�7�_Z��W"���x�D߁�,{=�H��?W|V�e��.'�=��y������YtuM\���/��r��Z�E�!�у��>�h�[�5��j3o�:ڋR�O"�l�uoZ���7��g&�rq¸!��|������Y�m����z��������omN7{Sk�r/�*T�r~�*+�J��?�~CW��������P�ʲo�Jw6�ɡԭGrzU�OH���/�M�h8����wL^�������V�^W��=�i�Q�g�q�7����h�՘EI���_��FN�L�^v}�J� ��%t ��a�aY�%-򦶬~��d4C�����x��5o��2Mϛ��Gf|V�M��������+�Z}|�}�����h���>��@��^�C���j���H/a�����<�#��S����m"S�)L�T��3�2O���A��;����rUUmЇ�*�F�/&�P��)TU��<n+:,���>�����Hj�1l��*>p�ĄD��ۚl=�q��2��K�-�y�E0���R�i�Hg ��>՞b�Y�ﶫ���iv��՝��\ѿ΄�Za��,#l >tt�g�̓�zXm�^����f�O����`O��z��A�R_o*�")Q��K��_VD`7�wO�����⎴��j����r�7|�Te��Ff�$�{�7E�X��s��I��ZuKҿ���Ę�.vb��T����:s���#W5[��ݔe�g�81�s������K�K�_�\�%$/jH�O��nΙf.��v�U+�N�����k_�,�]������U�k��/�c|VS|V}}��.�{v�rn�蚬zJ�f��5��԰��";�_	Z�>�H���n�b�<�;|*NӲ��1���@��L�RA�e�a���EjY6V	V�/:�G��*�"g�N���[�W����od��7�:���MI^`q��ԗo@��։M�5
km����2��0P̺
@�IZ0̶���>��l5A�U6����f�<g�8��t����M3s��ZԢ��6%ډ���ʜ���ֶf�����h-ee��/1���_K�vF�8�g����qڝY�p'�zWI5@� zR��eM�K>�T��P��t\��n�sz����%ܿ6����c���i���fO��q�������Ykn<I��@]��m���O�5u��A��Nrb�9��o�e�\t�Zm�x��u��Q!P��][bӃ��ٽ�\��2C��K��J�2;�./�	�f��+�,/[e�,[u���5k?�
��s�}6v$�|*�q��8��^jz�:��=��2���s���k���~�e_���yp�ҷ:��|�tb>�q'@?�NPp��-������T��h�	�g��K���y^P�D2F�}@p-�jOK��Fv������e��g�-]\U`��F��D8�<�1���z��v���u�̢hw^��M�B���:�i��y�-~/,B� ����L��Xޣ�~oc&:����q�s?ێ�q�h�8[ad�"�Cp
D#��x���d�H9�ʮ{�>W2�5���i���^��|
�/�
ְ8=��Kt�v�:rd߆O0|������W�:��#�AC� �tqG׿Q��g-"'[�����긵o�)����:y��S������ ��ܯ��������兼2��m�u�&B��D�$փ2F����!N&�qA����#�K�G����?V�j:���
�:��I�w�����Ȭ�b]0��>��M��??�̥����1��������R���c0ు���m�?����M8�8�ghlE�_�Ə�� AO��z��h�A���O���S�l�H�\��r���4�Cj�B�8�N�с�d\i��4��駔��&�RPo/e��t�XJH��Z,.��8�ԸË���SD7$v�L���X~&�8[N���s̛�#��s��p"�����8���<�FDD��Aj����g˼�saJ[_>�\8�Dj�Ճ�?~������������J$
���NV��w�?���*�(�äƛ7��;(p�?�'����]��W��]�4����U�p�Pp���^�^����ܿt����m]].�C��H�Qؚ��S�;���FH��.!�cpP�Р|)���t�
�gg�$]��K�Ŏ@�H�s@qʡ8�`	YW����5D���۝��ѕ��Α����B��N��O%��N.�445Uon�Ʋ�Щ�$4�������ǅv_��+.C�T�zA)6<��uu�5�ޢ��fU�]$��􋋋ٰ?SCH�� �+��P�/��W�9`��LS~!]���	P"p����k��-#=D�nz��ťW��5��� \܄�.�@6I�1��Z}�����Hc�2{2�WZW3��& � 1P	1J|�j�C�u[�;��@����]3�}��@��M`��o��ӝ�3M�D�C0�Ll��B�|����a��e3`��P�+�d�I��F�9����Sky�h�_�VG�J�b@�6���P|�0�Q9|�:a��]xZ�@H���}�7H���cmm�,BY=1�}o�9��ty�H$�;w���{+dI�Gi��m]������5��+���p^H��e��2b��쬬?DIm��-�t�=,j�f�J`6Ε�iݓ��b���\m����)+�����G�¿a�x��/��vBӄ�B��TPXHOj�V��=��ÇH)6���M����+ߺ�{��Sg�X*2��c:���jj��K�yS��Ǐ��_�jY���j1l�B4��n��ul�^�����4:������G
����}а��|�m�+?�]�?0���XtJ���3R���+��Gܿ)�hhj�K��(��3�3m�=@0i�jbb�+�A�O=Gy`�
�!��Qb\|�bG������O�<����
I�3}��
�"w�<�G�m�:l��>^��T��펙�|���&W��ɾXۏA[2��h4��RM�3^��\b�M�W��8�}����	��[�����<�Y/)$o0	��p�S�2�pLj(@F��$�l��Ҧ:v,���6��klj
��ӛoc����q�%C����BA�*���~On]x��YZ�~�f��i{���^�vs� ���h�&T�0�����w�=|��C�Q�iM�W��?2}�O2W�X^�G���������R?@�W�Y~5���Zd�PAMԑ���9�}?�h-�}cEk`������BC\{�Y���֩n]�A� ujr��Y�,oƴy�aIMZ�k
�Tq,{�P�	�+~+нl���l�(�����l�9��I��|$�w�@r9��m�_'�ꨧ3YW��<J���+����=]�}}��F���~�����a��	�\8z&&�ngN�N�)P3힚-���*�����ع����8�-�F-�빜Ej��6w�nі%�.
q^ӽ��������:����T �8f	�
[n�+���(���d<��m���K�����-�{X3f�82����T�[W��\�|��5�t��3�6���D5�_Yzz�������h�*�-5�8Ja��t%))I��Iz�W��o�ځ��{����S`d�>N�(U+M.��~|��U��Dr75y�P��!w�=G3�>6��Dl����}�cg$ �o;Ȭ�o}9[U�ƍ�-�#-��$�Mhp��:4�e{�	:7��'�(?��܄��%�E͊ڏ?��2�p�բ�<�9ML����F��^6��c"}|���RS^ZX�j��~A�b���J#F���l�qUS�O�mll4p~����� ua͕��s7��m���%����q�HY���3�ֿt瘛8����+X�>U��E״����g�j�A[��]䞣�[����y��`��V��H�C�i��A��#,F���z��W�,J�F�����Ề��:k��7n�8WfY�]�6}e{444t�������ޮ�q�aS�� �N/��.����ȷ�n��6��{l���3R�x�,h��u�P�Y����4��M�g��w���˿+��q��G"�^I����٘��c�^�)��f���A���P�R�hS�8��Ӈ�
�|1�ف�����1i�ò	6���=�Q��{�p�&���T���� +���F���l�L[��q��=w�v����ʰ֘�^^>�j8�=sʚ楯�oW�����~��`7���P���p.j�IF�(�<�z:�f��?TU�2^��K'+��<���e��Aq�����ZXI����{�(�~��_M���o��q�t�W"R�д�G��r���P�.)}� O���j	8��gce�WP0�X]Sc��\D�uez�&DI���fH�F��ٗQQ�e��|׆�Qt��?�c��8P���C�jum�H_6;7׾�H�ҥ���rM��R��!8���W��H��(�����ӞNߎU��)��*����O�	dڨϧ98n�G�Ke�`��1����� |X�F�yHH@�Vm$y����9pBd�o�)(!���s�y�x4��zxH�ٞ�C�)����"�	l헮W�����8͕X�i��c�U�%���(��h�9=��]������	�y*�6S�|d&�����A��A.���WD���?)�}�?��\'*����=�:�-wnR��ǟ�J����$>�= �v`���A@�+�)b��X䈷�wɫ��
7//�G�<||��zy����if���x��M�%,I3�b%����ͬE>Y%���Z��/(C��pۚ2
J�q�BWl�n��&�:�>a�Ɍe�i��9�}���� �r@���
����gzŁ��LR�VV�|��:LWA�*�v/�j0�+���Nc����8�o���r�S����qP�ִ��e�"��և~}�p�ɩ0�$�)�� V%�*)�
�+b�DV�HRt��	�g
��&�؁|$� .�E<��
pi�(�D3O7���..&�N6�X��<m�z^��׍vUi&�U��Sˬ���AQ���r���l�`��Fڗ@�O�
��,g���l2����
��9�*�j�IM`W�+�w#+���{��L43U��w7*�%��V�dYq���� 0���Y���p�豞�)�i11q#H��3���[W�2ɓxPR��s����S�{j�n��j�Ν����1W���	�q�	b�п{E��{�;�i�$���t3��[��Fku�Ť
N��H���٨`�uܸko���>�9E�)���A&�I,-�`
�z���r�>(��2�Eث
����rF�XܗZcx2E�cʛ_Y�� �6��5U�QZ΢�
����Z�,�:��p���i�p�:��$�W�����H�u�LYm/��1�4��+fH��6QP ���2�\[��hXP:ʛr��[f�&i�-�����*��Gq��.i�B���(Y��O-6K�x��{v�F���j
��]��g�Μy����4�7xFd���?((<о��z�ʝ�Ov�8=2����Y<�s��q��@�4s2��6~�+0;�Ñ��}JO�"��:��@a϶�5���er�.+�qG����\����é
\�������"��G4R�t��ߺJU\��Q����";'�7��]!		Ɛ��#"�7D�O �O�c6n3T��b�kmW�þ����ʩ�X��n��nsq��A����{Dr�YUa, (H!Ow�>`u�^����w�d(wA� G�{��;�Z[[i�͒ѮI4�^=+��Z+-�{`�.�;o�B��+�azh_�h6��jO�CQ77�z���_(4�ū��;7g����� �T�t8e�<H�]@��q�Cũ�����fgg6�/J�,jkk�w��1��ǯQJӃ�4�D>�7��eh���%b��o�h�RK���t����"[��E�VZf�R��CUu��c:S���ty�]�e6L�U��R�jM��`ߊ��ȈM��/4�Ȗy��V�W���%|	�e�)+�	F�L���E��E1M����Sy��l9ŵ�+ֿ8��8�b�%`���O��4E����^��������0���� ��:���͕(�U�^�ZO�.eRv���p���T8��#eU�r�aאpK�\a�3x�S���,�)�;4���$�:�ye�����i�#���߹����HQv�u[���~�����=�<|\��g�c�E�P��,���R$�4g��V.l���1����G��F��{�O� >J'}��W A8<�L�z6�Zr#�Y]�_��s-�4׿���������֜�?��J%G���{P��E[ME (�Z�G�Ib��c�^ށ}�,
К���ͷ�B��\�Ə�r� �fcc���oS���ވB����eC��� ���*��4Ѫ��+ߵ�Le#;lq�6P��48�HhӁ��i� �cy������Cp���h:���7�(W��?J �1�;V��Yafd��(jQ:�e��x[N@�,�k?����s5ˍ�pC��i!�w  �Y��tog�(�I���>lS���&����l��
����V����2K{����C
�_�x�m�4777����<q��ի�S}���Ĩ=�O��:�)Ж^�>�_&��)6�RSTV��-9O��y�}���|)��h'��4;�w�@�v�[3&�&&q��8��Lh�u1��-��-����n5)4��𭷀+=�/�*
N�j���:�Jԕ�L�#����5�B�_���n���N%����Eח��th�o���YҦ5AmM5�d�\�{B�E�kK��90�9��B'�&���#u���ᗫ��Wb�j���B�Cň��R�C��SU�w�.�'�d��M��TWWGv&3���f1M��$%�,.�QPQ���#3��^�Z�����R2^W$���o�|AEIa¬�v>VEC�b1��q^]�Y$\;p����Oh]9]��m����6��f׸����e��8&u|��H�9ݛ���y'7�#UF1��Zb�P?���a�����=w�Azjs]�J�ͪ}�n��e�%:ZQV-����:ʜ�cQ$�a�]7٨f�X����!�ta�Gh��lfJ���;�cVf�{�.��
򱕯:N;�ִ��ǉ�`���Դ�J�AL�u�̄nkC2i��Hh�[w{��H� ��D<s���n�s���չ���w�ٿ�s�\F�ž|�`�@�q}4*6��k/̀ei#����!�K�0��`�h�v$%$6�>x���0�e�#˽nRB��^Ʒ��ȐI�"�i�8��@:w�e����\z�<ϻM�#�v�`��+�����ߡ\�s%�J�VT|^��Y���\YZZ�V����XU�\�qD��ɌW(5�Su�y��	��BC��|p��[>VC�x����N��:���:1QzH����Cޑ�bA)���ߗ�m���d�qN��#�:h�����=yi�#� *,b�qo�]�B���n�S���'�Ѕ������|J؆)C{�_Ft��� �8��ɺٹ��?w�9腾�a��`�%�Ӗ��o�Ҥ_�QW�ENW^��b�gPC�)t �i�~�H����x�X0rmm�#S��W�,�VP���@���S�"�,i�� �X��K�Q��8�n܈<�_G�.��l{��V��J�I���Ev����
��;m�o�x_)�\��B�e��_���3b���נ�Os4��?;{J_�r�!��N�7�_�X����j�D��;�T�rF3+#��*u�CHfj����eي0���y'�>j(��3���g(ՔG�x.����*QRTʑ�s����"�a��H���Z�(�-�G���lT��Z�wq-�U<�%���b�����/i�\ G��`�����>z7D�t�`%�E����w��O�}}�c@�j�?�ܗ��{�i�|g�'�UG�dRKT�{�+B̏�өl�B<��6����9��y������sǊ �k=�@�5�2C���b�d�����rٗ��)����S�퀌=�>NN���7�d0����/aAĝꩩ�rgL��(pg�;��%ќz}J7A����o��V�y+s�`��[��B���������Z��Q�J3�Y� KY���3_f�E~_k�N�uԄ��^�$�n�(��V1��8�� ,�2��bp�������w�y@��+J(�9�T2�gjb��ȩ�嚯���@�%z*V�}�H�q��C�HSP())�7�N�d8�
��}�@�b�T���P\(wgY'����Z}Lg����;���w|_�+������C�6;?�q�?j���P�q��[T�	���&Ȃ�Z][�<�U�C���;&��^a<uVP A�q� �u�;&��B���m�X!5ԹW���E�1��~�HGg��Gw	VL��~��Z���|^^�$�s�Wy�����`�)��e�^k�C��H�B@:�|G B�\���l��q:@�uj%�w�w�--e�3�:�\�1%�w�w��tO�2V�b�Nþ�'�b� -�g��x5�"�9`����*�z���tck��a��۲EZ����H�\~A�	�ls������L�� ��GHx���]RXDď4ekck[Q�x�laZ8::�h~)q��b�@��H=��� x&�,8�����1���$E<I;��S3MK����:5݌9��Z<���鮾����,.˓�<,�W>T�ih��7
	��V�s�_V6f�j�BxhCz�n�bj���h]���KNƒ���Fl���i[pmJ��p~M͜�EU==�
�)(�a��g 8�Z����"��EG-
���d�֘��N�
p�윜��ME�C�/F���2S����+���)��yצū�7�|����uH5�-��KIm�-��!�]����za}k��<��V1�S;��6��r��Ba|�.e���o߶U-fv8l�4K��</�_�P�) ����]���#d��hJJJ�H.hN+��ut|�uu-�V�E-��82u#l���jzzt�5<���M�Q��Y,��7l�or��XR����cu��ϊ��P�{�
 'LĿ�8A���VZ0By�t�j1����y��������ԗ؞h�'��{Z�B�O�W����"�ʥ��8:9��&�A�t'ڦ�_�VZT@;�&�O�S����q+q��3��Y&h�Bu�u��08`s�k=��e�^�ٿf$�r�!hU�7o����TVAlZ��⌄�	ق� ���jRqFd��)Q֘���������׬�uR��dJ�/X�"3�QI�Cn�6t"m
�H���� $��q�S�אs�R:�_hNPT�a��Q/9GV�)P��J����/����8�ֈ}�:iNCM�6�r�JM�{sT��m�v~~���	�):�}'�}VRS=F���F��A�$�Du)��HSs�8��� ���[�z������&�/��10gN. c�]�����1?"�)3K�(U^�Q@x$^K]%	K�KjF���H�8y��@���ylՙя�pE�CȎ�O�l��T#Yt!d�d�~|�7��4�R?:#�y��ǐ�,v���X�aY�Yǒخ�ޒ^{N(�1L�w/'�"�g�������"���o����I����ooo#����B'F� ~�UgQ���	{�"���,���vG�]���%�&f����RX�d7e�%/���i�Gδ
�O,���Ǩ�H�����>��6�V�a0�)P��L�˿X� .vgx�u�6ۜܟ���l�����?PK   �dX����(w  +�  /   images/1485337c-0c33-4cbd-84c8-adffa1b45f33.png�|wPSo�.,�X�( �KT����t�C(�;(�Ho��;�)���Mi���йI�}�9ws�Ν��a�	�d�k�{�g=�Zk�PMu�kT�Tה^>ע��(HAqf����贂��/�߽�s��0T �;s��39
��)��r@ϴթ��@�c��~^�Sy�m�?H�����@����&%`������;��Ɩ����*.#9οdC6��񕭖Ĉ�P��?Y³�T��^Ե�y���ݑb�ћ���������.{�?ާ��<��7o$�'������������g���+S�*�%+���9v�G���4t,�
�I�@A8=(��#�2ڑ���,�����u-��k�E�Cps%�%]-
ϐ��G]����[�?ffL��#"�yd����gP�==���U�c��\�}�?u�IN�OIIy����2�\̗�GOWW�����k;�-�YϤm4b����}��Y*��h�+�e��/�tP�i.Ӕ�����#�϶H�N"�ii�H=�).�%Z����\��� ӿ�F���N���/� t����Z��N_�~���ӝ�hY�4<<:w��Gxx8D�J����ML����#O��	A��ҥXm��k+���|�*�[c1s�Qf�C	���e����~s��oZ�/	�ǥ��{����������rw�b�0�C�t#>#�����p�1��|1�8��;����Y��h]�/��2����$�i̍=��3$�{����7�����ܩݖ�%��}W<2��ɔ��І������q-ԕ�k����[-����5(���Μ���h)� �7H榤 ._�m*�T9!)���l5Fl��gR���

�_#�tw�}�Y��>=:�9��)�_O����`m�q�vM��R��S�t�8���������*g2N=�-ʔ˲↩�ު7��ˊk�g���\�j��W�7,%����L��ض��h��	�m��V���O�����_�،����^�,�7�uKK���Ʌo�pq���Ù�� �5=4�����jɩDs�!�Yݜ�Y���b���nx�����s�g[o�3�6
����?��g���;wq[�X�|�.a�Kn����{�>p����z����� ԧk�Jo4c���;���P&÷W��\`⾻a�[�)��b����FFӃN����?���Ó@TA�����]��!��%����v��^�����K�j<��/e���nSI��{��T�o��x�{�:u��7��_vb��,":��5���,v��VKN�ê������xZ~��s^{�z9U5)de/�	bQ���UmB�Tc��H����Y���{�Ԯ����,7����;�c�����:a�i�R��I�2�^�2Jq���)++K�P�ـA�MIv9U�@����E��#�6]��8��GHڝ�X��t�1�A�ڏhy۱�7�!��8�|�jiG��:_)�t��o55i5��� �*����G����cXO��[�W�_���+?nph���k핻:i��p���5dɆz��W�@qX�����|�c묋]��S3���Ɇ�4�W�<�����kj�nrg�}�h����_t�N�D�=�[15�Ҭi���cm�^��v5*ύXe����U�u���)���)�lPCP������Cz�w;W��d�/:��+۾O{�����5Y@r�,l��פ��7jK(^0��'�^wm�k��r�������_^F�z�R����1�`@�{��^��ט�����ǻ� V4}��K�6�����cSͬp@:E׆Q�Z9N80~�P�NO�����V�� ��;~���#<	��e@ɮ� =���zo�W��L�SE�2"j_;��g,�m�+��i��grg>2�ޣ�dF��1��O]�l���&^�H ڨ�S/E=|He�/"�}�X�"kTލ#�R����l�:,c�
/��"M����٤Y:s�I6?����!P�#�9���ˢ�tE�Z���cu�ZV�L����'u�f�R��״�el�y�}x��?������"����c�MjMgϳ]sHL��=ҪaNO�
7& ??n��`@��F��F���r����W�{6�G"�8�snSѾH�f��1��4�a��#�'�0�u����/�.::�Z��R��6�
g��=!s|5���t{��2��R>���M�VZ����>�� �M<���=d!�b���ʐ}�����Q�4�_W~(-m�	�C/=�}U,����u�����=����Ҩ8'
oz83�y�z����H@�ˢ/��;�ALɩ|}��n��y�wꍑ�xj8�[���u�H�{��;��7���ԡq(��]v���X��ʺ�c��٦�B�^.ݸ��o��dO,��Ua٩�2���}br�3B ���&D�h���������G&�=^Z�@�C�[�o>&u�g�:V�9�m|���Ewt��Q��҅�b@�m-�6��l����}���&$�p��=�zq�<�:w��+ ��������[��'٥�+BZ%����h����i?
�>��ɷʮN
S�`Я� 1ܿ�� ����cޢ克�=AS�d�"qz��3�h���͹����̷M�,���_�<^%L{��"��l�A�/,v�,��_���M�8�"�f�2m�V6:���*�����3�))Qz�{�`��%�!�A�;D���G��c�w.�{�9���csz�7�.W��Y���;��B��`��zMp*�H�;F������t�?�s,�C���-e�z�A++-P�3����7XĪ���~�l�F��g\}���"���î��Q�l�Ԙ�T�kǇW�h^�����y%��13>bZ������C@oݼ5�$�cr��ks3{�Փ(��Z��dֹ�]Ѽ7�������Qe@���:�� ��/n+���	�����jXD]vxU�^�&�00>�ѹj?��۱�n����"7�l^ٙ�-�� "����+G�ϩ$|q������%-�e�� r��6#�U\�����m�F)G�e�*۵��*�u�Tc��#Ϻk�Ӵ��&^�E�g/��I��-F)1�z�����ί���c�|���vl@�]񍹢���1��a�e\����i�F`՛%�R.Փ��DȞUo���R�k�e����v��I�e�7��:��C�=D���{�f|yV��TM��.��E+���<m�P�)I\G���aoh�K�������L�U�n��/��Z�|U�&�[C��&�C�8��yǠ�t��H�
I���WSfn<�)�^�v�?�e�6�ļ��ã#���-|��D�1�I�3E�y�����D�NI+O.e;6U浺n�/ ck��S�XEt� �Ҽ��Xla�cf#@̾%N"Qע�MR7��^~�Qa����1���c�ny��TM��`lTZO����z��f���G�jȈm�,j��Y�)<e!ȵ��:���jDt{�e95K(���Q��z|��N�\T #�#�פ�q��s�޿ٸ�����Q(��߭�ފ�k_���=}�k�l���JҎ��M�U�D@��r��c��nk����2&���o˽o��K���<��4�ٳ��� /Х���߷e@�0�"�2���4�<@�G�� ��ؓ�0���Uȣ���v�EǨ.a��~�-]-D��`�fAL8�������aUr^s�B���R�a1?vv��3;6���x"�P�]�o{��풴�%78v�En�(]�8�y|�l�FP	�nfE�ǡ&ʵ}2N.�C���M�&���N$
z��
wq^0u=$�-�*l6	�n�lj<�o\��]�������c��&<j0��c,A�a��p�cٓR���#@M������up�7�f��@U��,J�|��I&L�W�S#3��ha�~��p�|��H1�2��݊��OivV4�`�D)g��8#��w�����}  �V� ���T�ݑr��F0}�������p�eW���=�: *�QK^�.ϖ��l6�G���(f�g
i���#�U���uNq��
ڱ{�Ƚ�ЃW^PG�D"T+�s���������2pD3��@��c͋l�]���b��T*�����߻��.�2#���"MRO^�4�o��hQҘ��";�x��͛j<C�,-m��0����m�+��9{���-֍����4%�Ia���J���Ƭ��,[���_f�lG��D�n%pYC|���>3Yg<9�Ey->CgO����|$�7����R��B:����ˋ���l���D��aV֗�Lf���?�����hd��@G��}o���������|k.��Z�����Dd�a����1< ���#���[:^�]5��h
ɨ�"V�����#��h�ɶ�AFTl_��«HQl�}�i;��o�m��j��b�N�z���Ѧ���t�2]�ĥ��r#x�J�H��*�V�.�EŉJo��߯,�����
�O���~�:h�ie���+�Q�1�Q�O��W��x��>Q��Y�����+�t����h�n��כB���k���M��(`1�n��P|�z�P��4=��H�}����)�	N����0#�8ݫބeob;YSܪ�q�JZ�}�o�⫔2�z���-����K�
wﰆ��	(�Vy)1�b����j?��E�h�V�q�����b�^,6�[XtVĈn���]��/O�#W~��:&�'��Q��J�(��qI����������1�µ|�e,��B�,g��lQ����6X�~�r�:!o۵��]��Q�o���@s@~��jC��V�l���̛�g6���v��LO�n�9F�y����c-���k �R��ŀ���b���ٴ��'��˶��3������������6f�2氿h�7Q5�ÊMbY���]�3�����Z��Q&�O��K�-��<�=!�BӁ m}ؚ]�l�r�\Ṛc:���
�D}N���U�>�<Z=���Ũ\��o�0�t 
@n�o���l����X����w�,����
�CӿPqs����$�Y�"�r��m4�G�r�����~=��ب~8�n��DU�x���/2j�<6�Y�	�GG��H�f�|�\��̇��ՠ���0Ҽ�.6�m!�����l�^m�$��}�Ww�9h���a��J��@�$���뼴��l�C�J����d/��e�>3?^) x���M��%52k.��t�\����t���kS���W ��F��2���DpR��T��'�d�p�f���� �e���a�g�O�յ�*�y���*i�w �^�(!k���x�TQ˚��$�}�8�]�L���L�+�GN!�RR`�����pۯ�5��qOn�Ϟ!F���b��>7��i���xShl0~В��D�Ȫ"���iR���;���15"�þ�(�u��*F+7�#H��:��CI����eF>ܺ�Q��e2T:XJ㿪Ljy.D�h��ujyW���kϛz��DX��Wo@�Lϝ)\x�{z,�U�B�VV�Ȗ!��`)�0C����9��ii( ++������uƙ��t�Qȃ�_��I;�Qna��\H��/���A�O{�9aX��9��(>�F>~|9U��`���Pv��7fs�'�2�7���.2TW�s>��D���d&�	�U�+d�o�{�(F�p��&9�1z��G#�cuĽ�%Es�OJ�E	o *٠F�۽�5a����r°M�h�}6A�P	`ץO�,�������(��m�Bxc]'m���W ���!���݃=�wD���U���Rm.�U"�5�_����WꇷP�g���[�<�Y��	�jg��i��Jtn�t�,��#%TO�h�
��h�˗��H-����`�_�L>�a6��rR!ő�6��|�����d������
R�tC骗#/H,떾Y	��Yב�Y��k_B��U����ի�)>>]�
T�X�@n�G
V<�t�!1��E��1:�?
��H�W��/W�z��%�/��&.&eyW�%(�!��)с#������f�
J�-) �8���Q�S�E.*2{`ݘz�"Ea�{x�bQy�h��J�os�q�(U�4��|�X���1��&c�U|���V��f�p����kJ'�ۻ��������>��܌�n{M4�B-|,��������Ђ���*�_}R�N��wG��C�b�E��A�?��m.�(�:/�X#
�c��I��B'���+����cb���&1�%=���n����kt����.Uf�uT&ڑ�c9�i�Y�]�7����������p�;,�C��:���* ��m�a4���� h?�s�.9 [�j	ix�v�k�Te�y൷���mU��S�L�8^�,�VS��Y��ky!sا~��}ڨCߢ��5@����#����f��hj�1��������O1l���蠓��L z��ge�����Ή�Is���~�bp߱��|A�Ll�՜nk�י[���:��z�㥶#����B���'�ʨ.m�`!%�M\����a��W�<��:��rH({A����Bv�1(k��vo�GI�I�,��U/�U ���#���ILl����&YE+{�|
'�ᰱ����2�Z�?�I���/�j	o"�f�[;n�|���Oײ:���4���kX�Tt'��B�BǵTs�` י�I��r�u�W��X֦�J�ݖ�T��$=�T�,{���a�WT���5�'O��J�������\M_iY�9�}|���G�9=��M�\���hw�p��������զ�	B��4_�5��� ���N#r��'UoS�RP�b����!��cs/���m���T���G���zz����[�}�&g�v��c�P��Gc�e�C�y� 7e�t�<���!� ?~��5�q�>�zF���{P������h5ns�0��h�I@��ߝ��p�g  e�7��~[�U�,������F��#���j��0����ְp�2ouD:1p�o+�i�3zܰ�Bc�G�h��e+*�f$!_��Gv@��ъ����"�Y�:�O��﨨��|����3#�c���Q��{�Zll,�fny�	|Ks�	����+��&1�e�j���J=V����;�,F_�FLnBQ�"�{o_wԻ�y!���-)S��s1�|��39IMy`�n��G�$]IyT_w��Y���Ⱥ��H�hi%�7\�5�������i�u1��-+�,��Mx�1��`y<��*q�M����3#w���6�Bk�zm��A3��V�ۚ��-��Nn��W��|/�)9�Z�����C-�] :E�b0���S�Htq�G�ʽ�Ws��yTB=��J�Z�� �<D|�o�Wqp�Q�wo�Ņw�Fvk��BO$� �珎y��ER>��z��^n��=`6�W�\gU�ufZV��˅��g}�ɖ����W�����c�����isv����fdqQ� U�J��V�����t����ƫ
4Gp��Hy7�G��!��zX���0�Y�e��ڬ�	�̭&]�h�^wo��ʳAAy>�Y\�D��ڧ��=�?�6d�5�?s�E��&c!��F�u����ʝfա����{S�W�i�c�K��]�������j���kG�5�B�S�\}B�~���(�Ư:�[����%%��������6�5W��.]���5���먥��׮�W�����]�P�R�j��t�]��V�|Y8Zjx�~�F�x��A�?��F.�}s�o�5���<��⡫��K{���Q����f2�dO��f�O��)�M���X�Vs$7��|���QN% �)��d�@;����i�1c��2tD�6G��ԏ��s�z�j�ݺ�Ҿ\�y���(��Ħ�"�:Q�Q���3�^1��gy�^�vu8����E���?�%�Q ��D�29(�*��o���f��yJɣ�B���o�~���RT��0H_8���=n#F�NN0%��
D�x�ey�~���e%�V�T��;����tk�2����-��i��IhǣT5�7ۘ ���8Ul�4��؍-�é#8��Z㚄x���<.��C�S,�	�Y�[�r���X�W��I�9^�7 2�v�=�j�oθ\��w �s���򄋠z���$���`S���hIZ��}&�����'�i:�	_;�p�p�o��~�wQW R��}�[{���?��1��2B��Oq�&���PIk���ٛ� h+�9Yp��]m��{byΑJ��O1�c��ʼ�� ��w�VF��Ei�&��{�#���4�Qq�"uO�x*􅍾NG.�\��<��IR������*}_U��  �f���=/�N|�lF<3���O�Z,����s|���q���`nC��`EoU���C���I����P5X�/��K��6h��nhn�_�f����H}�ciO�����aCe���aM	E�Hk���l-	����"�ᾡ�-t�O�fc��Bc?�Y1�s���9����V����)T^b� �UVd�pS�o���ߘ��%����ZT�����qF>����6������-הS$�NIrق4�q�5��D^�6��B�R+��/��G���	�}u���r���X�P���V�C�� K��È�x'5.�KN]�F��_o���C�ɪ�<��SgڃT�X�&bY�n� /?�>�97�d>�ڶ9s�䌗/O3��&74�K�J��'�q uf�6�CO�I&NF��o�3d_/��E"��wxde��t'^�T�nD��&�^����|}���åo��W��_��1���Mf�z�y���ըX���$7E��������%^�i����I2C�>��04�2V���wa;� A$'#pA�1�%�n�%cz���...�t��<����x\���1�5/8vr���E�92>�t���.��y�~�{�,��)LO`�����JLT�ZKH�㱾�<v���!�J܀a��(x3w%��kz �ziZ��Z�u��s�B�JC��z��_bq]�3��=�5!$�(�;��#tx�z�n�q�D5�ʝ�J�#����>�/l��������$-kT�L�@Ña���)LhAQ��=x������|S�x�ɖ�%��)?~���{��A����T-�m�Y#y���$ӗk���ǍwD�8�Ŧ�	�	�j����<<�+�RV�&�ȒZ|�}z�fů��N��fa#��i�o�o��xab��z<ӌӹ|���W.z��l���Uq���к�!M0����	tyC�v���ZL�yo']�]?����2.�|�R��&7�V�����"�q=;�K������zy[˂��o����|�G��yǇ@r�1	���1�)�5��9
�� J��?��T���v�9�$�mNw����l�+Ýֻ��p"�)����0>��Q����a��qL��/��g(���y*H�(6��0d�>5
B��?�
u}%���i�a{���{0O��X�t$�R�P�|��;�m����ڕILO���Ui?}��H�tR��\�B�,Vc�+m0 �f�}���~�"c�&�M��a�\��8��t���\��.v�ޖ�Tvq'�ơ
n��8zv�w� t@;6�cO�p:v�l.�A�̼ݫ�|2�VL|�[Q��ή�<"�@�����P=�s�V�"�)����b֭���s-��:i	�2��.e�|��E��"W��̂i֯�׾��hy&��/�	h�2�U�>�X���d�z����a����XR���֘�,���;^���\��m!�WF���ޘ	�
���%q%�0r��tGm�
�V
�en8ޞ������o�J49�M���=�����-rl��k�U���<�	w:V8O�/�:ױKtq){��B.��_h	�s��܌�;^>�H�XM�	�o��IHS�)�4�M�'ϋ�U�{۳���ȃ	���'��, �=Ó���_�ZѺ�r�@R*:�"��K����Z����pX�ŏ�Z����؋�D��ߦ��2�ΔM�AьdC��m�]�vVl`�YMNw�I��z��P����dE0�}\��[��~>�Yz���$�ůӞ��{"<�ə)Ӆ�K��#~����^"DF�����7�+h��2�뭻�,k��wƟ��
����5�ϔ*�*���s�"�Z���X��l�ӑ�so�"PCv#�3�D����s�d�Ulr]���㿤)�7��N6�%YYOߜSIYvcv*V~(i�}��h��6~L9�M>q��9��b��G��4�>����3�)7��m���a�e��=^S�G������ix�qL=h�L�wN�8 y���i���e�
<�K-��K�lpn� ƯQHR���ML��8E|b�*a7�{݇�Gc)Q�	�ņ����$Q�9�09\ ٵZ\x}Cj�z�.6����ؤ>S��:|1f�����k���3*&��I��	�8}���7��ٰxSs�2�2���C�L��H�wwףb���0+#�Z�ۧ9a��+Z����o"��5�5*�"b������f=�B���~�F|{����UaF��[�)Ά����6�Ձ^��?�Y�?�oܖ��W�2��M~F��ZZ��a�e��ɝ%U�Id�x���~�"z�A��<�I�S��3mi?QFcNZ��E;2P��Y���j��JC�����f�)V!�O�Y����Xy�������N�i���$/}ל���l����7�댩���][�1!�y����Sߪ �03nlҜ1�6���09�V�L
xX��o�=�{\�����ڈd���s=r2d ;��q�Q$�y\n,�GS1�����S�F}�(�l�qT�ʗ����Q ��2�Z+��y�`MH	n�"ۙ�`K�O/�����8o���\�����S�V�/��{�U����.r�T�	9&�5�D�¯�݊'��[�D��
���j��>�IHX!���lS����5��L�8X��c�B�F���6���
��9wJ��=$ZDFX� 2�:����!�sW�m�9�o3>"���o�=���	�	Rm�5�Bu���"V!�G�ˬڡQa�T�B.���l�Ge�aɬC�P0��XF�o�ҩ�۫��q��L�۠�r�-��wQv�;�2���s(U���)��� A�y5�����p3�5Lڛ��\�~�c-mTB$�Z_@���p���p�����}�-������|F�jG���%�"�%���>��췦
�Z�g�=P^�LFu6j�Q��r���)��/� �3��U��G��XR_(���B.��ٕ��$2����<U��V��j��	ҭР�N�kl��}��5JF����ųU���0U&	�u��TǀQW��Ӥ8�=�d��Fנ�����ki	�mM��*AZ{�)�������e�r�LC��������Nny���	=����ņ��4_���Z]���dZ�����따ߖ+׋Y����PQU����<H-�+Ź�ǰ��ɻ�o�Z���ex[����������֪2��5 �/��SV�����{Ǒ*���)��pSJ"�xZ�٦<��6}�}�w�^
u�c�O���a��:>]fn�����A.ۨĦ�Q���ve"�םS���J�T����N2��dʹo�r ����5�b�I��	cT�!5�����3%UV����s�i\�\��:$�4�=iP1L����ã3,cEĲ1#"�ɳ����j�쥢�q�Q�}	�v,0���X�F��+������â�����@O�f���k�Q�2M�h&7]_� �O�k!Lq^���ĥzM�t� �����O�~0�Iʹ�ג\!����;>3C�A�Р�$r>�_'���U=���4����*��AU'o\�\)�`>�v8�U'�C{�=I�M˶�k�i��?��x!�O��F��,���Ϗ���L�&�����➢�9jUj��D!n�{�#��)?�;���rΗ��}���[q�*_n4��E�ˡ����{�����OTo ]�Tw<EK������!��I�Ï���U��w�E&`����U��/@�Nï.��n����5��!�&H����t{㑼�osX~k�c���9r�#���TF=L�A���O]�5����*�/Q��7ʈYŇܯp��0�B�����_�s�^k�J�+��%��w�tEʄG��=���+;�r�	l���F`������ve�Ʈ����{���梚=�-�r)�RLO6��2�?w�Cdh��e�-M���[�N�  �͵�P7��5*j����P�����<|w��."�T�?!�
��[�KBnB>��N3�"�D���(��_�S��~��y��8<�Պ�?���!�h"X1z�; ���f�\�TuEX=Ó5pzuGw!�N�$��]ɤZ����0��'km�!��Bm���O ���L��� 鎺���.��x-�u��%4忹(
C�.L�P��5�hJʓ��� ���a�F�Dݦ����!���,��:��_��v1��+���,_H��%��-�{#/�����I1:=���[�N������T����jkx�}�a����" k�r�u���/��/�"�G\���L7.���\O���
{���R3�jE6쳶}���S�c_�c�6��L$Iח�C�ܮU/�j&�x]qk�SH#6Rp��`��x&<�,���AN�I&���MM��V#Ҁ��v姱^����ɲ��
e�_�h�A�,`���b1���A��k��,���4��{�5� �	+ߞ��v�=ĜkhepY�>���^�ا�G0�P���/ז&���?�qŜL�0T�B�7�iv�9��k�����6��߾rח�:*\�,�,��
jh�xݦ�����9 ���d��Ŀ�H����Y�耓x2�&�ʅa�mKn�L��ϗrA�Qb�}5����ߦJ�r������8�W���U�w�ϯO�4��$��=���{�u�
hF.�ɜ��_�U�L�Z,2��g0�Oא�ڈ��tE�p��ڈ�����*|Ο�jS�םS(�����A;$[<��_ s���i��^���05*wl>�u��Ĕ�<����n�,����@�lb6n/E���ma'�m ���`�u�飽D�����kk�I�:����V1K�(�c�
�RH="�d���1��M�����Ot���]�⣵��Q}��I�=���-�lפZ_�0)��Sc����8���Iv6gG�G\v[�3���� �Tq>���x���c��Eg����7�U�dPҼ�'2>e�I��Ti�=��j��?O�"�H�OK��p(t����iD��D���΂N8�C����/{α�Po;
Yv�[eķ�a��������Bk�� !��0h �����sx��m�0�0c�y�c�fO���|�0�]�)>ZJtW?1�؟-O��wux<ҟ#���&E��P~��.?��2�Y.�U(yc�\.�����R<5�Σ������Q���s��xD_�0�T���Ym`�OE������fuy���}L��WF!���vN�q^��U�ׁ��%�$s��>xj��18��2� &��h�u�	����ohk���:l7ЯE(��̒�l�L�c��n����	T����'�������dS0s�Q�B@nr��s
�Ew��05�,�v���Gt2os스FИ�� K\���`kC��b�eP)+S��"�Hҝ'ͫS�Ȏ�<�%�h�y�Qn�ާ2��C�:�A�q�R�~��L�ƭ�4�<2���l׳�'���_A��2��XL�ɲ/�h�?U4uze�f�˶��6��v�q�y�<�r��q��ј@Bu2����_+���3ʤ���g䌳���t�Wj�|���&N83S����އ��DJ�W�sJG��\,��U���o�")�@2�~yU�K���ޑ�g $>��q�q8M/��d#q�u^c2�kS�3xX���"0h�(���343�(��J��
Wmܢ^zc��|�]�b�)Կ�+��%D�f��D�;�(����jY*��gm�,�[�U���m7�6|5��<]�5�]�ȷ}�������~�െ]JX���ր.:��f5o�F\�f�&�m,U^����f�gGނ�n<N��"5��R��D�W��19���U�#f�h�,.^!l	�p�Y*��Q~���S��X��4g�\���&x~7��o�ᵨ5��QcHuO���w_O@/���Y��� 9~szL�"ߞ#��L�~}��#c~L�X�/eז%2b�&w�&yM��7^��̘s��/{[:gE�io�O�#k$Zb��:Z<��}��	-�r�U�z�ח�|w�����p0�V^�IL=�rJ����?��ͱ��]g�I���&��%$���D���@��Z��fK�|�)	��a��`�O�0�`�t\�CGs�q$�����x����-=�m�}-}qY�~�^G�=Z�Z�]q�<.J	�j$"��\-?H� 2L`���p�����'ہ�=w���
@%�*�G��0���y�³�$ΰq�ּm���wB�����כ��醩M�_ۙ�=QG��� 0�lP�@�%�m>s�u���'��<� M(�?{n~6ߵ.�]��0_���aT�҇�_-R�ɾ�Fλ��l?�¨Fd^�;�uTZ'=��,����E�S����1<�o�D�������F7X�N�	k%kuz�!�^W�=�P�S��ϗO��(�2��� {}Y3:s�M����8��q��*��/��y�>�f����y�)��2��|yvq�)kJ?>��
���˹�ʿ-N=��餋|n7ļkH��u(�V(�{�α�.2�a�ٳ��Tf)ǽc ���ǖ�G�RdD��n}���^��{R鱧/@9�5�-x��[ A�4���(hC�Cb��D�<1�Gmɐ���)�T�����5*!�rci�������m���**�9�E����b���0B��n關��z7�Q��*KY��i'�s�]��!
#S�v��#������8�.��B�8]�h�MR����*���0���.r�ܔCAqz�Z���z��g�,[wY|g�(�U_��* dܸ���>���mcy.%V��+����?s���)�Ғ����0}��G��yO���E��\3V��zҦVZ7��f���V��}2����
��������u��.�
���HX�
��F<�t��|���BIm$6�t�"�?��Ms�:������W�G�3r��14��(g�kH�+��Wk^�*l��?�{��3��X���n�ct�y�ON>�O��EO��R�;Ғna!Mǐɍs���c1
��{JI�G���k�K�I���"�����~?Q�5���J�����e��'.ߤ��i�O��� �?92� ]����}���_�Sx]��0�#Ht����П��`���϶�^�5��[xL<i�yj)cu�p�L���݈j0]���j;$�����w�?(��|�]aSl�ȣ�Ba7���ԧ'���3��`'���V�j�Y��c�*y"��qw3��+�������ޮBA��ŅBt_i9hF3g�תʄ�	%_I�?�����<,���[ە�0ბ %�E^l&�}�ph�J���2�YG������^�<ˣeL&R�_k�o���c9��vC���f��x���LBZ;���D<7�J�ߏT[�6�Gm���8T��T�����R(�h��G�7><,����䄻�ў�mg?�@%n�4�zL�Ov���D.v%�~�4og�w��6�.2G�p�B��uS����1�T;��������ӜY�ڸ��5�X��Q
��^�d�)���x7n�K����(�Бi̬�/����L�m��yBɍt� ��&�� �;���d�%�VӚDq���O�Ϣ�}�ISk��K�JH>�]B��U-��!��٭�&>�1O�Q���.�����CC	��C�	X��D�f�EG��� B��87z�V��W�D��x��9p�a��rӇ�2�9N����6�����Oψ����|`r?�x���+C
T�S3}d�{�����3�8ZZ&?s�q��"��u���{���g9OTym񘛸����2�I@65,��^��[R�]n���Z�'��;��u���b��qد�����8� �
�aL��L��g��̱�o����{�����[�<U�"�B���/l����	}��_Iy\�?�{�;_�����--A�Z�u����yb�m��0M\ ��p�^���	�4�vDv�{Sڲ�n�xLs�8`�qS�UR����T��Q��̟�U,h�7�Θ�̹[O?�Z�Z��3(�"fwoDm�����xǡ�m�h����X�a�8OS�	?�����K'���;�|t{�gp�e���c�uXW���)��l�z��p����I�}\�1�=k�uʤ�04���m��%�
�*u��1q+UE�s�'p�^Wn=�������`/��fEl���xuE_��,E��w�`�4n�2_�4g�>���P�ڥDg��i��R]�*nT����o"+�u�f����H��@��ل�Z���F��v5�v�H���1sB�Q�1��V}s��Қ�׵㭹z5^����\�#k��e���ȩ@��}8�f�I�"fF���������+�[�n_�;},�`�����KEj�O 4z�*<���X�A���झ�ݝ{��ÂO ��F�KaOY>3���>��5����QBb���AQj^����ޣn����l�z����L`N;��U�KĢ�k�
���Ku��RT�g�)͏�!��i޾�sT�O'��#��G#����i
O��7�@5�N[�)�v���=���On5{n&N��R�}Pי��=&A�7�ϭ���#�H�|�f�N�I&@�T�����
7��D���fĴ�_)G���w���������jrk����9r�RP�IWQ�HD�(�!���L�  ]�=jh�A�H-!t1�B�y8缳������o֚�<���.�u������PQ�
7g��D�������B�_g��j[��qB���!�5y�/�g�U�P�˃��[4�����Y����ṯ��F�X3D�����n��e*V��l���!�<<'C}�fg%� ����� p� �P��^�B)j�?��\��\������|����n�{чK�Ȑ����x�Jն*$������rG��̢z�8�Qmk�{�9vj�sY��k�Վ}����o��U�Ϲ`1/��<�Fv�W�cY���ܹ�������>~���e<W�~�`�^=�U=�W�D�M�;3���*� �x��K_��C�4������uӧ(�6o�zf29�6֎膿�� �9��M�z`�!#�9�������}B՚��,C���Q���c��)|c���}ҫ�g��U�Q�9^C]/R�U�������s�ŎUx��r���pG�A�������w��ß�~g��vLTF�y���5²!��-6�b���1���x�&p\�I�{�^�_x�?��t돤�҅H��H��~�wl�|vU>�9�k���xB����e�'4<���7vҵ|3ɸs_���w|��W�#�UM�l��Jl��Q�	��wi��x�u?�L<Z���6�'���"�Lx�D��Q�`KˇO�!,�X�>h}_��LC�j�ّ�֑Y�$(��!���t�"*��_��SPyֹ3���f�.���;əp@LWfݪ��0p7�u��撥�Wf�Y�aN��X�]܀V�F�4,9�?�
�.�d{����&����i���Q�M�U܄M ���Ym>�W?����9�Ӵ�k]��u�7�J�0��"'~$X��t��K�V}�JR���]b�2�3��Jd:g���r���k�d]��Ĕ�ڎ�wͽ�k��n@��b_���w �W��×1 p������M�������GL� ����t@-���{j|!���e�\�8�48�����Քj�<�/,Y�K��r�̖tz$�H4���L�����M�+`"�����S;�4����ؤ���4٩8�k�&����ڈ`����@6���3����s��[WDl�ȝ3l���t�8�o&��Lt��Pa羥Z˕A�H��N:u���\ bS����v�͎�>����ۏr�U2��R%o���d�b��czS�U�ě1�L����b�r*u���c� ��%�q�!
�٬AGB4YU�t�4�RZMw�j	ݻ�"G?��2|�����Z��XblǺܝ|���I�-�9������8��ae���m�^D�=�q�a9{�/'x$6t��5��Лte5\���o�!g�[ف����Gt�ֵ¯0�g�h�o���ܙ1�;[���{!9a��y7��+E�/�eG��, [U�V6y&�J�Mc�eOՐ}̋��Y!2GBE��^&�]u�m�a�7 �/��]�5��8���m�4�� ���������e￤���a���c)�Y	
�O��du��S �΍KI�uA)�y�P���^��S�VqZ���l[�&�:�j��T�,�$���5IH���9p���g��me�r�]aW�y���Qq�͝R�U/��T��|_���q��\?�'y�VZTl�,)*q���.�����yK0F�����`4�I�@~�s<�
���2Z���Um���0!ſ8����!Yo_��"��`OQ��D��g��h��.�4R.1~�t�ė1V��nݕP}�9z��)xI'�"GĨ��"h5��Ǩ@�[�z��$�d5`�Ĝ~��ͫX����ʇ١�������S�A��6��&��}�}z��A8ܣ�D1˛����q� �M�S�ZFV��ؾ��%�b%��6:+7��`�o��Z �	�.�y�U!~��D�ݵz_�������7�8�Q�����]m�ryq�e���gu+�	 (d\�F��u������K�����ɵD�m�S�6y$���I�Y����P�6`��}ӷ�k=�c����]�/|���Td*�"8�}�I���*/��,[�"l�槅3����o�",c��#m(��l0��(ON��C5���ww-�}�{�ez{(��wX.1���	\��LXU""�#�oʇ��x���b����W> �/wa+r�K�4b�ןD�m��:J���MP�m������7�Gه��N��T��#e=C���Z)��&_4jX/�Y��3�l�z��r����V��E?�~&���y-R
������)�q�
�0*`j~��/�q��LZ����&4Mp&��gi�n��!M���/�"�l�[̺2�ݷc�)?��P+�q����h�S������j&�o��{l��ec:,��ߔX�����AK�6���rG[�?Lq^P@��m�Ȅ��ލlEo�fb޸�)hi��ƪ�7�ݚ��gn�Z) yHk�_������X�E��_���s{ a_%�T`׳W5?Z}.�C;xD�x����^��ʀ���8�!�CV=~j��EJ�]Aw;����~�]�F�����>�vq�1� HEHY%V5�z�P혡�Y�|�^}?PӍ5ISpU���ѵ�6E_j]��͚���-
�Pu�u=1�3�m@Ц�WWn-Mx|��"�7_��y��ј�DU6���N�Ho�m�����q�>�Y�c�6�ޒ�t���w��4�1�K��f��zӸ���@˴�۩2�?��@im�Sj����Yr��c�D��T�by8�(��?��q�:�!�˾��42��TSҔ8�cI{�P0k����_� �M�H�
�g7l%Q��jw��:Y[�.<%�j��"kSd,%�6D\F��S��h���e5�}k	���3�i����S��HA����fϰ9àt�y㣭��"�89���:kn_;)k�s�<�紷O�(nbV!�̖�*�E�"� *����i�6O���o��D��4H<�.N�޹��ؠ.��e�N˵�F1J�1O.�_�U& 2)Fc��(�бґ�1 ��3��fF���$���d�������gJl �t�h�/ݴ�O�,sPvz�'/{�������U�ݠ�H��A8��P���8���)K�{��i8i��Ȃ��6s�AZ�u�#X�7����J-Q�Ɨ{U~���v'!z�n ����I���*B�i� y _�&)�G��/U��cs}�S�∴o4�5	,�R�\!}Z ��^��u�����h�I��X������h��4��H���gW�on'9�GHH�+gv�"S��J�{��l?�YM]�]	��&ܱ����������#�:�r���:�e��R�P*�zU���5��OV�g���jZ] ��F[�rFv�7�,���-��KM����%��5 �
���K~_��ji��F��F�q�jW~�c��G#r�q�g��%�e��A������`�i�
�s�]�`X�t~������ss� �q')�*�j�~z�,%%S%��^5���.5�+�`}+����V�~�G��vXJ����L�$2<)��k�>�t�2�����ͥ\i�#4|z�^<R�8*�n��l��]�U�1,�l���Q�̠{Òr�Gkבw���u�
a��b����R4��̪�.��8�*�h�7���L����q@���G>��ןt�a�W���9�'�oC�E{F	Hx2��:���_���RH�rW�j����Z���O>V�\
�q��_�=�.x��*{=?��0����[W��5�9���H:N�BR�1�ɪ�j�cb�+�y A��t�9���U
 0Y?Z��h���m� o_���� қkv�����GK��1�ha�3Ո�jK�������u]�e��s���y�t��Lx��(���ˏ�,D�rܪ,O'?>�si �3UE5�&���~G8��a5��4�ޠG�Gq�:���˶V՜��Դ�G�����'S����X�����2`T��^6��~���=qK;}���Yg�u���3T-UM+��9h��|e����n���A���|-��m�;�Í�����9��l�M�����x��ԟF�h�r�M��/�p!�19?�^)*��b?�(.
8{����U���<5|+��x���덵�I�VX��@����dSz�����ኀx���A�j1�z. (`�>X~_E>e5cI$֋b]�b9MՑD��n9l>��� �t��AQ���r�W��	��o��.%�k���]�m��ț��Q$��������<����w�e]|K�Ҋ&e�՟�^}}���5�,F�rUHVm6>g�8�ԑ �t_�U�[�H��5|��6F�5�I�p@�y�/�ʗ0��G����8G��n6/U�FW���S�&(	��1 �YTX��L�ϝ7� ����1n�Yt�A����#f�p.q���;!��AiOȀ��ٷ>�,�5�s�5WxT�Z+?�=�B2�R��:�؝)u��o�}�)�;��z�-�/caN�]��� ��(a��]�Q7��5�%�2�8|��Qz���<�SvV%�:Xp/wk^�4�XwE[��!5�O�>}23��,�.�;����/��!���\o��hm`�Q��)����uN�u,�d�GެdH���|T񷃇7�`A.�������4)@�}�ʣ���G	�K	a�ϼ��r�9�8-*
����{Du9~2�{����L8��}�H
>?��t�ݣ?���������C�$1;��t�cS��@��puiO��B,�f���D��YP�-�aIY��xJ�5)^.S6�Z�8�S��;��^;��t"�<�M]��"Fȗ@��A+mΨ�_��9��5z+}�����˾�c/��:�w��D�e��r��-�䉷���{8@�}�ٓ�fT�LͭbZA9���	s-�Vl@���I3:Py�����w���Uu�HGX:��ݤD�T���j�@��k�Ҧ�ܠ����Z���C�9�vD�Ļ�S�=8W|����<��J�p������gN������~���M�^4
Z��j�4J4Xo�����f�7F��߭�;�8������	p��&ݪ�Uό��Z ?-��[�i2�=0�d����#:@:L`������&iӤ�O"�nk�$��+�gm;����0(\�I	[{;����2L�9�b0b��<3wm�Xm��	���8��� `��1���8���z���F��i�MjYH5�G��j=��J�7",����-,�ļ�ӌji�%�,!n��XTc����F��ru� zg�*Lb�#Ζ:+��!g�W3%bVu{�T/�d�/:�S���Y�E@��
�.4�����mJ�iI�Y� f��
^��+�6ؖх֛�b��]Z���$�(��n���(���ͫ^nZ���\�G���=��ńU|�l�{�`յ�}�"��̞�gV�8�{�k/�8��6�02���y-�$�'�a�V|.#5��֥�[u�q�%�FP��d�^�y��q�;�Q�0��?&��D_
8��'~��Z#qc!f`|U��&rasƀ��BC��K�'�ۚ��f��N�Y���4�Go��7��Ü�k�o����p@w	���6��ix�nwF�i�ـ�Z ��Htf�>�I����ގʻb%�����
��9�%�#����ez��I�u򨆋]��}  iK��6q�y�4R�Y[���հ�<�����1l`���8�-��!v���I�����CG�v�҈\]���|-��f��am����o�B��
��]��,˻w�W��՚���M�r7(4����-	Q�_>ӡֹ����GNq��;�T�����w�����T�;1�!��Fak���4��L4��U��m�H:���.b?���-��fK�3<{sĮ)�>p���^��'.j��xwb���
��k�á\�i��[�
�|
u��qaW�H�B��q�t�m��Etx�pdk��ڼ�X�h^�u��	��#�x����QK|��J]t}Q�l��a���=�^w�_����J����C*;� ��[�3>d�k���p:�c�W�E�Q��ǋ^z9&���T�nHF�u$�(�)xk����ҫ��������UO��pY�.�����o0��%C��{+�p��n�TV���7��l�Í!?1�$�׎�ey>T�S&�7Y�>�%o_&_d�K=�z��S��Q�y>$f���kw�9��}41�A"G#�1����:�4J��z��烏��������gyM��� ���8'�l�r���e��<�N�>?FI��2��
��/|3<3����TZ���p�Ƞ��B�2"�Mػ�X�3�љ��Y�h�?'ez�kpa��� �bgA+Ymj=�6��^=�O ����.�k�??z��F�-���0SY[�jg�}��ѥ�gU�����&�P�+�~�Z�Dv@��=���K}Pc�B�����Ŗ��{mˤ���O�7h�	���f7�3 |���V�(�O��%���˛N���=�����~!�B>�)�,����4�!-d-�rc3�Aߥ���)��r���_Ы��Xg�}p�˷W�EFE!�_�����<`��^#PVu8�<��T������i��3�4�9���Zqŋ���L�9�vHi�!Þ���Ĳ	�<^jC�4
�9S���Ɇ`�����7���@�߿�����j׌�CCr��w��B�q���+�}�Ϻ2��<	,��)[�⡲Gk����k��s�XD��J��X�\���P��"�w��k��pD�/�uE����?TR�ȇ�߷�{~��p�	8`N��� �o�b�ƍ����u���]�jG�z��v@P�][�~���`�B����%v�`��+�x����t^5�k{c�ng�e��k�$��4V[���K��I.o�<�	���(J���.�/�IA�b�΍��e��,޲��t��Q["��\��?�b�'�{��4JD:���&}�vr/�V$��l�i��4/����OZ���}q�k�l��[2�	-�%$�1�w�6`���uo��
��g�q�- ��ȁu�KM�үF�k7���3Gk���O�MT�h�p+��?���?Q�D-ts9�5�'v$�s�;�dἥ��>uc��߄�G�H����O��q��Y��.v$z17�'���E�/Yug!���
f�`i?���bop��[��9"Uoc�GWp���}��ڢ6,�Pw���ٵ3�(�.~#���݈/�o��V�����2l=ve��I���x�4+���9�M�?}�ґMoZj��|�Y���+�� -�Z��n@ ?���q�^oC�b9VUzf��\������������B =t����b�S~Z�yqFƓy�������ϑu���O�:�O�Q&Q�<~}�?4ĩwڄ�zo�/_��O��|ރGm���͑�ʏ�C,�����ٛ��܉�^��ޠ��g/]zP� � �㠂���_�;Q퉒R�ݮ���R�	{��Kμ9�q[�Yx[�/�W�����Aq���+�o��4��;5}��222	�����յIxg������6K��GQ��q�3M=ٓkfY��^m��\�x��F�\���䵽y%��J����,Ǳ�����,Q6ɵ>��E��<���E1���|&�p"���|22WE�8�8�ۤ޲^y�x��K�|�m�t��Ƃ:3CR�<����������"���JC�P��pxc��aj�<{d�*���#��0*�s(8��u��y:M� I���mK��=o*�Z ���0��v����&1�m��6
��K�4�������
D�y�T2���n6?��Og���;h���\�����%�0�leصk�g�|ʎC q38,W�<�y��]�~���:'{�pE& J�� wB$=��(�������)vw�g�̌U ��^�2�+q8q� j��G�o��c���W]ʱ��gv!M��;��W�(�x��Z�L94����y�Ov�E9���'�׋���w݇��J�����B����A�-X� ��iɑJ�֝X���c�nk1;�-]����㋡	n��B���E_/�!��Ԟn�Ihf�M.	 � �>(�ݕHP<Lq��͐���7|c�s���"�����U�o]�^���$� ���3=n5�L�`��#��+�oTX���E�%)��P4NV�%{[.�o�=��'�6�oE��R#vC��C"�\���0JS�8�K���
�O��f�y`Hy�����^��&n�g�_癮��IՋ��y�(.z��\6*���Lz	��=��m�2<@&�9? ���51�i�ݔ�k�6�1��Z '�脮�M���.�<��i���47�a[���5�<�C�9حI�ەh�3�� �� +9C ��۫=Q�0{?���&��3I�V��[��#8��g�@6��*6�Z�'2Zqۋ��	11`�}��i/?m�^���Gv�̍���{����0f�U��-���f*:�(�Hr,ȇ��ùb�,��L�P9p��Rpu�/"���L\�έ۷ۜ;'_�@o�@��{��fl$/"E�t��~�^7��*`#�J
_���Ͼ��P�G�e�l.D/�~I��މ���<Wp��M���I��eO2,�ee":��ζ�v"$w��J8c��!K��Ke�!��?	�g���E�Ԭ�@�>��w�R�su��)�פ��\��&%K���~�[��+KA���l o:���k^ `�,:�(�JP��`��{�X�t�w�9�7G:��(AZ��l���[kY>Һ�Uqq�1%D�����_�����i���
�.C���׼���Y�&W��B�:|� A�X�4m�:us:=pqC�8+G�^��t�y�s�7F5������m@9o���۹g�z~�kgkx�Yu�ʽ�ۍ7Ϭ�I){�Q\5��r�ح�}���4SM�^���;�e����E���fi���f8�z?�	��=Z�D<z���YJ�s�����໒,@��7/��UD���+ N�{V�]��r����/}Ț�Id#��?o�ޓ�s]��O�u��V��:���@�*��S��	�,=��f�G"����p�p���˃�X���"����=EM��~�/C��~8J�����Fk�u3�#��x�3Tl�DP�w���"ӅW��s��pĭ�ij�^5��%b?�/��1v��C	)0�ƒ3|[ůP���#�&��.aC;���;��s�k�3��m[#PƐ�Ə��UٯV�>�ǘ?�d���/̣�2�u���1��[^'�>����`|��^��-���v5Z�k>�3��>�����'&�2�b5g���3��c�)m�Dq� ��W�ϫ�kl|���6��-С^֍��[w
kIA��|�`1R't�#8z���H>�#��o�Z3vL�����7�BXz5�1���ꍲ|��hH��o��i
P/��wN��������3cf�����T�o���
�?۬�5?�t�)V�1*d->��
�g����z?:�59!��N�>�{�k�۟o�`�O*�|:�
@>���K���_�������/RJ(���h����@.����ɡ��6V���G[���(P�����t ���^����h�|�������e�/�5��Ĝ��*{]����/�돏,p��c�N����BZ�S�k����'vDT�Xy~�I*��v�晀@;�H�MR�t}U��'&"-L#�����(!} ,vy�q���Q� �q��h��g�X�N�ȉ�j�C_��n����Z���*e�G����g_���O�\Їz��>P
�R�Kw���|D��ˣ�j&@L���V��;�4� �� �+^|�J��+��$9KGwA�F[�����H�y��m]�1M:v�p4��zg���̗6���@�㒳{ ��*^�H�,;hr����7톮�?9��!`�nI��<��sl0B�CL��̴�2�xDO��'(H��=�A�۫�dZCD�]�ؕ0��3!����N ��
��9�d^���`�� !ngJ�㈊��<� ��ѝ�A����t��F=�k�I;Ӣ*�&��ՅL�D�ѫTi�<[vo�I�w�lk\<����}4�b%� B�ϢA>�}>]>��ي໨਌z`d�f)"0����͹g-���I�:_�9=
��}���^kF%}��~�E}����CXp�п'5�@��\�(<k�n�D(h��<F����a���E�
	���|N趨%�8���& :{�A��G�o��FN���BYYd�^,>ܑL�j�w-� �VV�uacy��|/Lb���3!�95��4Z���>�������,o �kK�8���$�vS��a�9<U�����ĉ#&�����*�o���TE�QU���(��{�pGV�돇bm�*,%wg�ʛϚ�������M�]�"��O3�{�TUZ�����i��n_"�֭�a��$px8�O��]-�.���3��C���\�N	�����w�}(��^������x���&=��5Bp4<��ic�!a�#�]S�Z*4t�L�Ƭ+���kJ�xf��­�@��Y7�o�����iQHb�~�%t�M&�Ĉt&�܁�LD�}��>Nm�p���ަ�����Z@�I\���׬r��ol�>�l5|�_�D����^�|>���Ϥ��P�K6:<�>XTF�ȶ��蠖i��W�M��r%l�����]� |�wV�߈����Wb?��35�&���.�7�7n�~�S���de���
��_��If��i?z�p�R��~1h}?��T�`���TO.ع=������W<Zh?d�7��s�)�����k+������dfߛDf���d�h�8��
�zZ����u7i1���/�F��c��v;�Ҟ�b�/k� g���[��xK���b��L$���MwX�1�#>��ZZ*��cb	%�'v�)l/ ������B�\�� 4���i�0KÖ�K���V=9*>��ox��6C�.�$-F��E�h>�M֚�%����	��#=ާ�F����P����{&��-:RcDSρ䕼Z�K���XK�`.�n{TU�w���p��^Auo�eCC��5�,b-�q�?GGN�̴��:�n�~���� /�Z���p7����'��8R����(Bt�=��m:��-��8G�(c~��ΧP��+3Ϻ�'�1.���ބ�'��=d4���!��sTܶ�q@���NsJ�/ο��g^.������(� �49pQ�>l@Eb�n�;�O�GT�bw�n��2VѸ�ʤ�K݅��큄=�{�p�����.aъV���d�`�4��0 �j������N�Z��~�pʃ;иZ�nv>����_��' � s�:����� ��y99m�=n�1'�"5S�ܓ��k,��k�h�������}t=Gg5����\�ݔH�}��ڥ���C�Ҕ��*�5w[J�~��n�����v�^����S=�0�'�����dA�Yh���^�i�� ��M�2�M�隋�y��g����U��l+��V�$v�^���*b��5�~�Z�7̻��a��~�ޅ�|X�i�j�>3�����Ȓ�冧{r��ε�&��#$�`�A��s𨜐�!H�T:�uRv�RnU�LPS�]�"�=�PqH�Q�,�Š�7p�M�:�W*\���P #o���Ѱsd�o�!����N^��h������Oȇy�/4���Qe�qp�(��Vo:�d���oH���&[�����U������W���c�LU��Fm�혟8=��(��;o�5�	j2�ʩ�{1��~{)�l6g~E*���C�������K�9u����f�&��mmU׀��{F3�n�"M�$vVZ��! ����=�|+�n�O��Ζ*-�U`���`����j%�$]O�{��r�R�$m�EORC����|$p�Jw�����ɞ*������ZC��D���m�Js�֗��Nm�j�>����äT�	H���Bp$S|��+�VZ�Qx�BI4�ɶ�AHX���*�^�7Q%O�Ы��͙<y6���*����i�յ:f��^<����z��0a���P�īU@;��O]���ҍ����������M;_��-���s �؝�>�'��U�=a�S!)��Dr�`Ee��c��qg��!�ى�x#}��E�#�Q�g��:��&�w�>/�}���W r�U�����s���>F����w��O�m[��]%|����k�A5>R$7dmm5��o��� �`d�ut:1p�JNM'��c;x4��1n�6s����vG�ٯ��9�d4Pw����಍�9���uO=��+�.���?�?�&��z��&�Sw������">qh�}RRd]�IsJ�e�*�PQ�k����e����Q��ܑ�ͫ��嶽u��/N4�Y�f>I����]�'��3FsF�4([M�އY΋�����ʂz�rrڑKkkT�:%Q�;^ȫ�d����؆��ѣ�a�U�l�O�8:��𶢚��S���r�5�Н`K�p�Z\�NE�=��PG��w�D�2�I�nfb���vp����p43���Zެ����&���oM�Y�v?^����d`��h�g���/���(U�nU#�:�O�[�+8al�&�����׫�M8�������ƞ��/T�m�� b�]���'��o;Ѷ�	���-Z��D���S+e#_><�t���u¢J�6#/p�zV(8Y7+~�oS4��}��]Vu�3�d̵)�VTTx���v�������j:��Od�V�;ۛ��!��n Q��.f�uߓ���}��}��Ķm��5Bz:��̲��L����rh�!�:����"R�O9E8\��t$2�~ Ҹ2��Ϳn	���ZG��7�����b�:rX�G��PJ��!	��;ã�oQ��g�z��]�* �?�&��%L}+y����[�w�D�u(�Rϭ��z;�L/�o|6�`xhb1g�\�|5l��|��}��ݶ6䤼(� $������^����v?M�3��Dv�+��g�����g#��%W<�� PK   �dX��@� �S /   images/15a77ed7-bb2d-43f5-af73-2cbf4ea4040d.png4{<����EfB�[V�2�����!{�l��;{DF�k�B�&��+;][\{��?����<������|=�����p�����(��,������ܺ���(�!x���?xO�w�o#��/�_#<�ݬ!����vN�pKsk^g7��M�;�]���3/����ߴn&�6< S�ng�"����R�;��QQ��*A��6.?6?.�.�2�+�o̑k���|z��b�R���^��fs��A�m ψ��k��ذu~�W'�sjX���,8	�}�����������	�U��D�X�voQ?xc<�-���6���h���	Mrļ���Ű#��j�l�%%�HXKJ�/��I�`kU0C�w��W��o:w�9��n��5�+�ᡋy�z:Z�t��%��C &2u��:>�zk��X"�Ou �w��Z�j� �.=z�/����ھ&G2�YD�F��?}y�n)y�C��*v^qH2���ffo+g�-���h	v0�+A�psۼj�X0L��ϑRS=S>|`z'w�S{!�1�7IJ(���g��Tq��k�@*�gee������x&3
��W��H)�.����2>�I��@�m��X��)u�u�����%����CΤ�U�1Ҧ0�����(�*]]]˞�	=]݃+Z��-�Z���,_�Sb�����{�����
��٧���5�Sj�C���1����t��J�4y�D!�ۻK��P���	�����:�ދ����f�D��>���=���X[/�u�moU6Q�%���}"f���	=���<r466��t+m������Q����s��`�H?��=W	Ǫ�����%(��������RQg����s�桺_Cy�����<�)M&q������!��*E�M�e�_߇4�ױ˒��>|(VJz�����jC-CD8M0+��<�4rS7�,p>][[�1���?�mf˦4&!�:�=0[�~,^�r'>#����v�S56VW�(++�T{q+��׈��ODHH7�q
��z$���3�}��Sydz�2!�Fk[i�}����*�恪(���H�T���<υ�v���NEd<��ZHil�k����-�P�D�JG�D6Χ$Z���XI9V��Wʻ���J#���Lt��:I�I��Tx[�wQ,S�NOO�����;2�cX��B5P���.Z��`��t��<ճ$Ol^��,a���.KB���3��
���Je��UrP^B�X�(~p�,���g���S+���<D��)��-�j藘�/��GN����`��"G��.4��ׄ�����%(�>�_��sG���zC&!���k[[�/9h_���L�zJR\��N5�d�̦���N��C������������-�� �kes3`�xg�I��y�avY��=ӕ��6V�F��l�㩔8�C,���LRL�iO�H����@�sȌ>�vww�Jiq���74Ĝ�����
(!�]�49t>���>:88�TA8�		yL�)JJ�;ڍ�r��珎�>Z�V&J���?���a(�,�
��P~0D���﷕U0l�z�{�pJ47-٭B��õ���Άm�ʠ:��p������>ݣ�� %�M��ᒳq�m��zIX+�SX��#��!A{��=~,=49ٌ/����u싁���7�߬Qt��Q����[ZZ,0�i��h�T<�$�i7Q�gUs<�.����u��S��6�$;��o7��a� �-��2i��<^���$|* �u]�S]UU%�����1.g�{3��MG+��s)�C�zx��
┆����J$��8��`��oví� yc�m�$�9~b�h����8�7p���Wׅ�
&�o�	��ԙ�͠kHy��{\��}9J0;�_�m�嵵R!�����kb�j��W�h.G�H��g6��k��,)���m�!�y`��?u�3�1>�L�s�a!˥_iYO��|7 �̾�<%���]@���B�R��i3���S�O�`(if���L ;��?'+0��̶+�w��R-%��*�J^���[�n��Ih&F3�i%8�m��[��.�c��8�w��)]Iz���4�@&m��ol���[F�Y�-� ��S�R�?�Sm���)��	*d�)Z�c�Ǩd.���"���5�J�5���dHh2I!�+��� r�!Ĕ��Z�8e{(H���I��+.��� tY���̠5f��� �� �)�2(),\"�QTG��{���ijdѯ���BA�W\Q!-i�F8MT-�@�o�{�|�T�Es$��E���t.Z\��]�nܸa����v�1I�lN5��z�*E��3  �[$ע��\��@$v4�!��d�m���eq�����]���e�YX�v��i!u&1�i���%�3�|E�+��Q�Ϡ���,{�A���j�:��k�=�Z�HYE%��]��
lJ��7��b+�xy9ù��)L���ͭ2���y�2���7�����&@#,��;�"��Cs�P��%~z���*:
��������==5nf�$��3\�v��v]:�s��_3'��Z0�6�u�{(�v��vd~,���?�-)���{����3�1e4�_���T���]:��XO&��<I����ږ4��p�BЗ�;�l�Z�ɉX��V�!������+ŗ����`3�φ�vQ|Wc4�;� ���=z��#[y$��r��9�/�zDe�݀u!�T����fZ�5tc�������ޚ��Vyb��ӳ�s��k[BF�E��p֩�R	���
�}��1�1QmR��?B4SRR����=/u���"|Bq�W\�U_8�~o�a���=OOO�#)�!.���:���R� 3�0�A�s�5�X�U�H�(��"��y����#	Q�9���\�^��6��k_qa���k&E�%��xnNf�/0�xi���A������˃:e�V���}-e5����ԑ�T �AT2��L��/kmm��U��k~tK�hg�}m� *(Xt���}B��.��eUҎgS��^#� �u5��nG�Sُq⃰}���ޠ�?�ˬ(��g�����vaO�IHԿ���vO�޹s�Q���䗍�^����%�q�p_������R&W���r�:^r�G5�$�8ɭ�n���~	pN@�?o��ƳH_��@��%O�%�rW4�f�+ěp�_�e,��r����K��v���1�pH�B/�����{���o��7���	�J�����_���v�io�u�a�{��/���R}0GX��B��*�h�k\Ei~~���sE�>@ʦd���BK_�IK
��������8���`���Be%�c����,�9|E�&�=��f?���˫��rC�$�	)|����KKQo��D222Ԇ��i��=�q<����gz���_����me·�͌[�||Qh�4ջ�؍�5k�+�/ �~1�|�F����9�������""�O�&�.����0:CYoF��g6��������g� �N���� �?�AV��)��4�*�6�\J��o/-�^��y~/a{���K�kt��ҕ)��}�4�����*���T�? s���}����] n�JУ���Sy%��ܬ;���Eq���쳅���Bsh+���=�Z�A�U͜��>�� w5!�N �D�ٔ"��:���n@�-���%%���r�R��y�\w4F��m�go
F��� �?��� �h����m.�S�d�<��Z��,:x�j��\7�^?�Q7c"p~�ȳ�}��t�ӝ��~��̒�*����&ǿ#����d��{���GH��Q������Z�E(���}{*��"�o��cf�X%�)����bnK�|1�V�}xyqv ��vc*���G�bv�?@�
�dA����$@�,�x��PĲ������UOz��g�7�t�}�g?n�i��^���{�A�r�k��5��s�8=pE1�Ϥ�WW�U�6s?T�-����r�ρ��(Z��z׊H4>�2��_[\�"E��$�e�Ԓ
�6���ؚ6��kbb2���6Ue��4h���󛻞�(�mQ���N�X� g%KJ�?��^�bE%sےc�
�H�0���A+~W��>��H����@�h���{&��׻�D��zJ������fWR��\T���"~S��zK��ߏ�җe2X�X�zN��5�Z@KC
M����{Q�hh5��#���[CɢGkm��~��%�Ѵ�V���zC��H^��@�紁���p�';5��=NB?���.A���A/`p���^4d�z�7��W�=n���*�<T�.*��x�^h7Q�xz�Ħ4�荅=td�}����L����Y26%-ի��( K�s�do���o�[F<��W���;�ԻZf�x>�u�0ͷ���4���#	��<�DĘ�Âd��O�;��¾*ͮǜ�gf0\�3{��q���!H�8%$����o;n�4�B%V�9 �~^^�L��]"�����'(��a=1G����[:���y� Hz����I���Rb�O�
��'e�h�?�v(�+%jp���*���'P�����מ���e�op�=��.cŝk�9d�b���L�����Q�Tc���>+}S���}?)Ӭ>�ri ��j_:y<g���4�5����=��3�Ȧe8��~|��\RR\R��̹�9t��)k]Lw��hl���-��z���k3<t1�8 �w�^��%��	�v�"��ie���(ɲ�c�Zc��7��	���Ub�u�7����DP����l�ΘC
e;��]X�9�t�]o(�X�Z_00c<�=�_��N�u&�44�ռ�Kaa�Շ,
�ڭjǌ_H�ׯ���/�v�]����*I2{��g�ًbQ0�� ��M\ 6.��8E��?:bⵔ�j�7M����p�P�8h���Z,)y��D�bK1��n��C���y�>L�����6�.x�����d��Z�C*�u�>����'G��TTPy3�K�gh2	�;F���w}||�ka��Y�я�˛�~𳸫��Hr��=(9Q��$��u��]̓{�~���̾�/^k������j����|��V�ze���e�3�V_d�V-3�d!�ر%�U@�w�䶽ٷ�8~k�猦��������[&�.����m�1��G �7fڮ"�uJ�t�,E9���B�~'��<u�Ԝ���h�l{0��C�<xPS�!=�y2mLw����1�e�?�O��p���Qa���^���o�� �v��W������I��`]��.�'�9_�������,����-�� T����.��:����&ӵ��/�FG�\4�����蚼x���&<��j{�k�f&�9w*
H���{O��ʏ��,�@��x��ۤ�X��T���^$����hx�������~�pj�A~��8���Θ����c�h���1G55�l�L������69p,�Ƥ�Z�u��w�e�Tn߃Q�@��ܠ=�NQJ�B9��~W}��#�ۺ3_��ܒ'M����:�Y��$��x.�,�bV��V�@Mkڊ�"�r)_�����3�H�K�lTz��0��\�pV�l���=�h8T����OO�RE�4����%�cY	 ����h}b�ŢJ�ItsbߧeW�?o;r]7��a`q�}Y��r�k�彴�K20ќ	�~��V#�v��TD��dm1*��0��H����M���Ԉ�x����ɧ��Ҋ�- �� -����+�YC�C6��u�\W�X��E���	��\�9|�,���٨g��^>kgy����5���F��bza���j�#߻��{�����-�rzz�A1����x���<��g���u3����=���� J���]WzR�U�ܼ/�\���c��s�]0.�ѥ�9�-Q �GrX�vN�M:��'-3Bl�I��&
<)�z���[�Z*@�/�]�I�E�K�N0HJ�F`e:`��'>�'@�R*'��ђ} ��r�q܊�� �@
�}��+��0V���߭�;��*NMN�s.���������(���
�q�w��t����m��m�yY0
+�v�̓���,����B:b��$�6����S�`�<~b<�W
�.>����yא��W5\�l�7����p��2�!��
�Y*�@��܉/��v����+N��,J���e7�,è/�c9�Ն�o<��2i��/,|n��,؞���
�e[KK�e Qo4,򦁶0Y�4Ո��B�2���/..�Sjf�����w��CU�E����t����Ө��X�	p�j9��LN6� �$<�����Ց��7쭻?�C�xr:���n�����'zK���1�G�K?4	�!f�ٰ�ci��OpX9�#E7 �s̀E�0�Ò���٥/5���|��xs/A�U�zP*�1�����
�ji���3g�z�s�s���(A���hV���*EА�{�r�E�=��}>�Mn��I�5�t�4h;"l����G�r�\o����;���� ��f&���l|0eK��Q,Ю��ߑ�.���SBj�ӆO���h�u]�>[wϊ��$�f�1�i@����?V�Z������dbb�  �&�m��E�!�9�bF{.C�_���M)���c�*E��>�P�ǡ�c����F���R�W�*��g�^���@�g9�A�������3�,	ўx��o����t�ò��=<^����q�KT�M`Wr�{&�cmm=��/i�u�
6�..*�V��eT���1�4s|3��Ŭ{��tL�f K8�1�@�p�n�kh�D��pQG�;�Df���PJn�m]�_f,���X�K[�n�+SDPJcc?�[R�:�� ֛kjF���E�*Q�����2SD(%=kU�"����؁�A��b��ْ�j�,�{;<�UP�h+L-\�:�|�6>��%a���;+�a\�C\��������a�����ё�ҦbPiҁR���a��zS����s6��7��˶ �wqk�#c|�nS=!�{�yZ<�gG��$�-=*=�}���s2�M�
�;���B��936�|P1N���{E---�`����0NMe0�(��eζ�GD]�^@"�Y�|�R�֭[�m�.f��m̜�<�Lp
*{�qv��A�$G��?�o��[me�\M9-�	7�jdjG4�R9�9gAb��v�~i�&A��W܂�'<���Χ-TM˛F��T��B��t�%;/��ZR8����z�� 5}IK{�Y<M�y@S̔�W��!訮6��iT��fD��ԫ~��Z +ilJ�0T�u�շ��y���@�ra'y�� ��{Wd��9�!�V�[\�P��v㔰���ן�Ǿ�����T�3<���Hd߫M��F��LoV���ES�~�a����XI�.F�w����w�Тe����H��X\�(9bNveN1��=$��N̰�8����u��G�ɈB�������?��s�.�y�ߎ�"s�S˿]����e���~�t���RR�v�Ix�fm`5^n�]��Õ��������N�i!��n)*��_f�KG��zO�=^{��L]�C&c�^H(�E��B�tS!;�`6��l�Z�s.��F.ތX�fk��m�illlMT}�0�Z�ԟA���f�y$f�
6��[/��p��'m�3����X!�ָ��PO��A�����ò�Ӄ5�(4�|N��}��?/q���C)s�F#א�:K�G��nuݵ2H��=1���3:�#�:-�I�mn���`�g�p�&� )�0Іʓ��WI��&�<���j�~*-E�X�����ϙ0��8�{������b���#(�NY_M]�}h��N�� �=e4ZK9�`=����v�mg��;�NE��F� ���Zj,Ƕ�����h5�]mg06�x8�z拍ɆR^۳NҞ�.s�O--"=�rG�0��@ ��g.��g=��
�s�%4���v�,h��?�<DK�N�IX�l
�59h_�
+��6jܒOPz.�����1��Z}Rs���@G[W�:6M= ����vܪz⊃��&��9�a�85(�����2^tru�?V`���7�v�C���pn	Byh�j�Hj O2ywyc���{M�a��|�2��QR����O��Q&�!�����Qʢ�i�}�DනN�G��/~R٣�O�>���(����In���2?<�&pI/3�S�@,�����C��d��?ONO�c=��7�:�VV��(;@�=&�Y��@u��L�kV?h�늨�A��eÞ��[@��re�Mb[y+�������s��������)��+B�bZ����y�����}���=��a����}K�6���n��sTWd�(ꋑ��)p�gG�`u4�ҲW���{������@���ճ�d�ŧ�QoHN�Ζ�m�KJ~���;u�|�6 bUI�Tn��U��ê">V���,�9Q�ƿ���I�(�ԙ<�^�ZG�>�.�ƳĢ��	r��o��c��0�Éq'��b�|��i�l����� s�F��'Z�� ]4�z����:r���I��[�]T.�(s��T���ڍU_"�!Z2y��J�X*)�)�Jp4�����"�2k�#+r�JT��l��#�=FO�׼-3�wTN^��j�Q���<M��C�����L��d�!����\`��B;�.�ݾ�<�t��8���2c�����*�56od�tD�7h����+��kA�� uz��Z�	PDupp�i�bX��e�W�l�~�|��!�`�\k��ު=Z[[-PIwK*jh�>�yǰ�7Z0�5 JG�%7X�KZ��#R�@�Q"e-��8{�^Ӣ�(Gm���4"D[��� �2��m@�Fq��������� v���*�ٸ�bm]��i4!5��ؗ�W+`�Z��Tt�`�7�˴9h?;y a� �+�yY'C'v��19�Rj�% �a�e�2#=7�<�ڀy��1h�a
�[xo]�J����=�q�{����,ۺ��4&��΃Cbm���$<�[�����Ռl�>ي���_���4Ќc����g'�-�:zz��|�b�7�g�|�ı����s��]^o���}'���\����>l����#�%o*�UJA�-�����ȽL����lP�P5�l56�$9,�WWwE��m���.�;�I��\v�$�В�s�+�{�Ғ�9%lk��<�&�����'�i`���0���^׌�]�pQ~�.�v��#��������\B���O���B��T��į�ۂ>{+����7����V�Ļ����6(7�u�1E���r�����r7��k�~B�7Њ�������VC�ԓT���H=�� 
�t�K�I/��tr�.JV����\q;��r�w�(s��a��C�2cW�L3P>ܼ
eee�K��"�+++�m�p�7�٢�y>���7mp�A���;ʃbf�r�zJ��n\)��N[D�Js�s~�ȱ�'j�=Q���`4�n�R)�-���k��M��)����G�]����?���M�ާ�+%��c�A#pDWjz�e�o�*o\-�%�aM���NNN�#(��Ps�\��'� �w�PDt�{���i����/�ɰ:C�k��+AXCT}`S���fd)�1�f�}�9���W �^�4��5~W�i\��~Ŗ�t��vf��������:Z�5��G������8.	O�7̀�M}�#��INtJ���fZd�u����f��2�*��!k
���q���Mu���B8j�1<���n}
�)wo?��)�#z��kXU�|4�Q�e������I�w��#�BE�{e&-]���b�'�B�\�|]��蚅���"�v����Ⅲ�7�L�n��~YT~d�_���zx��������7��Ҭ��O9��Vf;B(�V�R�҅�;����׃ëO�c��@ՔD�<,Q7�\][+;Xvػ����A��oY�p)l����븓c�Q���	3+�kz��/����w��:w�?�y͖�H�I�����+��&��Ʊ��\�YK"� �C����?m�m�YJ-���!��q�:��R/R�����Q�x߁LS�`mp��@B�� �����pN^>����'~R((\-A}��L`�;v���D�����>�}G�9�I���T��) �ə�e_;�6�LKZ�\�`��#3��u�ra���M~�$����!S��F@��ʻ���x����j9�*Ql�&��m˔eX���(w� (�Y&I���<"��95�n���w�T��bŔ��������n|]�U.s2
��������ˌ���PqUIf��!�x�0D�x
�_��lj޹B�X����'Jɶ��l]T�t�"��H4�K������������-�����#�T���m�����xf8ޜ�j;����^Wɚ��4U�)Y����b�#Q<eX`�p��H���� ���Z���>QN�o~k�aC��|�z�h�xg��5p�yp����Yaa�,�j\�W��Gm�����ڍoFK���1?��W`���$���F6���,��<��{k�g��;���c�;A�S�r5���_��3g?��Y:�	�5k (���*�3��@�徱����M�1Q��������Zy�PyU�v�jI)cu�Uz�ߡ�*%��~ט�%(����� ���������߇���q�[�g�r�0�ҟ��IA$W��<�1��F7�t�������o�8�����J����|..v�E�D�K��A�<ۻ���Ƚ�P*�[��U%���V/3���b��c�@����8���5C���8�ĉl(���8�&]��W5otE)�^��44,5
8Y��Ht_�ǝi��i+]w��gc�#��А���,u���\p�%
 $.��p����g{���6+Z��.�@&r�!A(�"%%%�*j+�WV�@]i2J�y���>"3>�+�B��]�M���7r�M�nb���$����8�9�7�O,��Xw`-���=>rĘ��=������"�!��V4)Cr�#����w9�mU���b�t�3��:��ÿKKK�L��UU�v}��q��B9�L��d#(@�ɻG�L�����}����vg����ʸ���w���lP,\9�Zx0�D6���7�k�������s�<��W�Qu�eg(��^O�ހ���y�q��#g��h�.�ڰ���l�D3��n��Ʊ���Z�����R<O�c�?�����X"ދb)�)t���].G���I�,Yڥ7�7�(3��1���@��͌�"|f������?LD�j� b�ym��6���R@�� �9Z#��/;�����'�R��߿�����|�h;����HP������j�X�#6��H[+t_d=��$y��ڍ�Zq�a]]�GQX�x�vq ���7��kr��aE�A�����2袃������c@�1=~@#?66��{�i�]l�I3�K��k+(�^<������)��/#[R2�Vd�N�=T��e�B�>��Q6ꄩm�gw�HR�]�L�]f�K�G��･E9<Qk,:��c��=��Lz�y�W{�ˣߣƼ&Reg��F�".kk�Ξ~R�u�NM9zzz�xMz��*����m�7^�)��ST�����e�V]����
P���(%Z������iM�X-�~��8ʷ?�`�)�ɞ�!��W�⿣�rwj+���`�.s���i]�}�3,N�J���:O��͎H���x�F�W]�(moo�h�oOm� Մk�oM��I��TT�<�?�O�]���~�Cڋ%b~�?�����eS� ���v�Pr8:��S2���U%��}�AU���\��D���e�����yg���������p�A	맂�Egy��w���ގ>C6�^�Nf���R��p��Bg�:R��7t۲��n|sy�kcS������6���Q�����h��|cH�z�r}VJ�������D�9M�9���Xh���w��qF(��*3ID)k�M�kfS��[�hp n�(sW'�,�ko�0}��N| L�#���?��v[$�S�6UW�nn�.��[c�ĤL�Am�4������E����r���NR
8�LW�%����DY&ס����+�&�ٔ��V��f�P^Z�8�3G���(9?�]�a��@<dSe��߾����ԧ�)���gȫ_��&��M������z�����^�L�x��7[��W� y���0F
�o�����0T�ތ/�!����z�zsHQ����-�}tsD0�����_��,,��G�GK^uP���ov�A!��a��)|��n�����2�<�t���a�P���6Ye�::䍶��^0�����u�>�L�3�gX��Y�C�3�	V�;��Vf
T���x��d��8�7����s<��:v�G���~�G>B7X���B�V#i���2��Rpwm�Žw�ݶ�cF-�J�1���y��#�K�|�#��1�?bepn����O�L�����T۹����-��XЫD Wb�M�s�ǎ����.���2�n�9�1�c���ISY��B�`/.�����40�� Q�r�im9�ח �jƯ���`�����;^f�3 ����s�'��RK�{#ޏY�6��
&j%�Y�8bZ�q{	�CB7�qDSk�v�9wt�E$�\ϛE>�Ԫu�rc��j0�}�AKVhwǉ�a��N�~~�s�:�ط���3�EN�1�F�9�<�����a][�Jc�v�b����hؼ_�:R�r6A��h��A���������)���lCО�&�o�;̮�h�4�{>:���XO�k�^�]\\��������yAm��_����b�̀�y����	;)`Y�Dֺ���#�����hY�2�a.�5L��v����g'J�>�įEZB�X%&l6�n�~R����f�+��H*����y]�?�X��-�A��Q)��=o���S�M����<A1FÃb����NҐ�Rפ* B�=O�n�F �s�n���2�M	(�t������D�C�GL��t?ct#���B���(5ӵ��Q4W��p8�D�j�ۨ]����?�{��3�A�}��oaa=WDЉ>^ω�
*Hj�up���Ȝ�:��y�_��wx��Շѩ�� idH*��p羅�]S)//�ȃ#o$Ì����tAc��ְ�B$���_��DC������ҩ�Sls�T&J#ț��~�N9P�ʐ 鎘8�Cկ����" [*���b�����.H��_��[Y�Ki���������/~�g<6��aI�_�m�b�6:D|�Ѧ�#�ע��r�L�D���`Y̡qޣ�:��5SJP#e���~rW|w�zF#�}u���x�K��料���޸t4�����s���P���6��S�<vVR�:~`@����Nt/� mԙͥ55�F媈��4�𗺺�1�9�b����EU5��5����	���%dH.?ó�6��9#�i�^�UxN��j߈7U@m�6��}�r���9���.�"RK�]6���p1O����mX A�[�J(���|z .ww�>�lV�|��F�N8��mL�6@"�z9��F}��F��}��n���)/������A���NG+��-c	��LLLqƿ��.���i�&1}[t��D�9��j�X��A'b�W�T������K#�9+���`�'vqL�%�~=Cu�_�����|�`p��b��E2��Ca7���5�,�M_��/b�?�b�ib���c!�+���������$nj����w���D�#&/r��Ľ�zC��l�����'��yxʜȶ�v+�w	����Cڇ��#o�i����Z��b �3�A��|�/����J��k\\��MPG�S�'iI�Tا��d6�H`J��q
�o���DϢ@����2֫P:�'��ͩ��&ϭ10D&��_( �c ���>�(���&�[��� R�7\�|LC-�����~����(��4���v��Y1���;;�o��J���qQ���]"W�[ S+�!�5���.���7���@&����&��)6q���r���n�`����gM���1�_�`jȥ���Y͠-�AN�,�P��k2?�ˑ�O�,�SXԒ����+59f��"�N��h^f�u�����h�"���9������k�L���O*0f�q;U3'��r=		W(O�\ϲσ�^�%�������n�*�E�2լI���?�h�	n�����y��U���Ԍ�m6`5�� �p��
S�#V��A�#d�|=��3��b�
�A���v#C�rݻ�"Hޕ3x$�Ayb��c�6�K���!w����m�a�-r�gg6�b�Q��|/EL�,h<d܄!�{,��925��#l����l�z2��[�v���'w�$E��u8��6���p�V����cP��]��l�x�q�3�耂1���t��9���߯���R���櫔�����Ū	��s<�(�0'�g�&��s��$������bݶ��/J�¯�2����rO;{�&�q�ޚT������q�Զ���'���V=�+�P�d&A ;�'=���.y��gl߁Z�0�]�"�֬��P͖2�&ӊ4ݘn1�v�G��W�ʛ�][�ule|��N��y�6�,gA���:�bc9���m�����ə>�g`�Lf�C8	3n�{�"R���4
q�H���y ��{�/`�	]���Pe"�,~���F�6n�^��<��)��u^��?�w<�ֈ�7+��[��h����8F�&�.�i�b�c`���L~�� �+��8���,��e 7ا,ا�篴G���� `��7Głb
�WTD���u.��W�b+G��?��}w�?0^똯��h�Ŋ^�ML���ܒg.Tۛ~�ܼ>=8�oa~�ȶI�������2ر��vP�(�.�Eo����.�{Pbv�>==�6j��w]H���H-8�Ro]OϺ�#'X$������m᩼��A���+�[�Z�Uˌ���h�0|t;^=���㦋���s������F����t�Nޝ ����8��1�b�h������j��^!0���U��Q��	�~��hyKK^�LIE��h�q��Q �Њ����M�����3 �Oqo됰&�ĦTC���Q�D��2��!�b��l��A�P�5�:%&��G���*��|�@�Kz�CM��s �E<;4sL�v�K�0�B���	O�g��uVT%��g�P����ҵ�X��~c`a73Ps����X���!�?٨�=6'W����N����#�^ӥ�~�tM��<v"L��B9�^����
h!�Iц����Iz��5��_�����y�t���6�k ,/H��t�`L%]��k�k�Y�Cg'ł"��>�P7�&���U��gg�6�`�ߕD��i�K�o����6���ټGq+%BgZ�bi�e3ߡ�>���"n\��d�L�Q�L�X���zz��^㞕�q܂SO�zk�(%��P�5(�����pH�\]���تrĸ�P���]y��:/�Nul�[c3�����K�⃤@�@A�MO,49&j7&�d�JZ�3�Yp�:����r�M&�}�yF���Ǘ������'\��w�:645��p������D��4��@m�O@�1��+^3R��ŀ(so�)����g�G�h��P_Sߍ�<��eG��+�(}*��.���IDNNG����Bk[�{��?<@">b�8�1' 	*om5!��b�}Q�������&�H6=��Ţ���a��fwpw�=�
1C�����fyk�sR]�j�S�9^n\�h�Z����ϑ�e���w�εe~��zʮ�����{����X{���������:��&Y[��'�@|^�3�ŉ!�R=Ѝ��&��&��.^�*b�:��J{���!'��\��誗E�Pq�y�@ܫ��ee�]|%OSc�d!A�`2=�+#�;�xh!�߬����������eA����>[���q��ʌ�ϣ4�ya��p9��� ���A�Z��lJY�g��cW����;~�y"SY5�^Rn2���+�m..&m�B�Ƈ�_\�P��a�h�e��;���4{�QQW�gQ��(O���)rzz�[�F�X��ptt0��b@	���B�����U""<�2H9p��q��ŏh���uF�{���ْ�Z�~Oo�t�>0FA\��-F��g�Rr�l<ԙs���6��f���SQ���w������||�W���^�CF	k�������O�ñ
e��%%T����X��7 �#) �GGmK+㴕WWW%�s��[�/@�F��k��ƭ�	Z��
�� ;�;B}7��Gߚ�C:�8ql��j������a��^$w����c^�%�8	؀�����_�z{��dr�͜C$k�CU�m��n�AΣ��cА���"��e�~�E���
��lS h���lӀ�<�lQ��@>9Z�f�"�
����c�,��\�~��mjj�	b�!�gs}�Aľ8@�A{��W�Bh��C�#d��'���	8D4i����k�vxn�k4���v�zaw-���.zlqޣcR����ޅT74��2S11����n�����������xi-�n��Ԗ�,R~�L{�g �F[��F��Y�}o���[��K)&ޫ(�F�}���+� o���`�s����/(:������sƔˍq�Zo�/$�<F�ª`�4�|�vG�"k�����lme�w��2�$�=�l=��],��A��ip 3r/���@�,�n��j�������f��Q𩰰'i��AR%���v�|!���P<�4�t[T��T�R@��	S�\я���rmcc����Ma#
b�lB�Uaz����@n[[ ��`S��#I��cPU0�� .�ho1���{�oL�z��d98c�{��rZ� h�f�2RL��,*tD��hq��:K����*������`Z؞�a����&��-��u/��%`.
���?�66~�9	ąP���`Zl�&��������'�	�~"m�1 ������Ǒ����b=� !s�x-u;�6x[���7Аc��Ώ]��9e �cobF�>zj��������3S�Ɲ�v��8�,D����4���{�@��a�� �W�Mm	ĭ��ɓ'4bظ��ޗ�CՇ�Ad�B��&Ki!����ۘB�udi0�'Yƚ$��U�,�}�dJk��Sa�-��3������^�^ݷs��s-��}��q�:��iN�B�L,���VW��e�ya2��n/ 1�Ng��������ӀdK��j�ٳac�F�U@nV1����ߪ��`��.��/�g�G+p[t~:�Qw����l������d���~�A5���t@����j�/^h]#���rA��x�I�V�hh��[�P\���.�2�/�vg0]j}e����q&�j�����"����!,�P@Ό�z�tarQC�a:�=����}����qz��������O۝|��,�
�#�H k�/t�M��P��i�i=�8�S�V����@�Mc
��2r�:5��ps_+����5H3��A�n$��z?�汣��/\�<tkn�
WS�,F�?��:�W��7��m�BC�Y�P�*�(v���I$K�}�;��}�h�rX�?�|SO2o��y���17�O|xD#Є�le�Y��p3��<�t^Ŵ3�us~pm���ş[VO�ԭ�"l��/���Wn��u=|1�Q�IpL�iֲ#\2��^ޮԺ�}�G}����nz���P*�m��ķ0��2����1&���sn�f"�S���	Ց_�hR&�4^L/���� �
z�=9�IY��R]M-�Hb���w�&��J���1y|��[-�1�٥d�	�}D/�"ju�h���dW�n3<|"x�pO^Ҍ��Z/%�s�2Ĉ=��,�w+�y �lB_���y����/��-&T*���pa#OkR<eR�}�������~OЄ�R��b����n��QwQ6�#G0啋��L���|ͨ��h�~)9����{t�����=�G��8+"�N�CB��_Hv��Y���ewvv�����V�Ld��zO+�%%����^}P��d���� �'L����V57�����+����V����1����2��*۽����Ѓ~��x��KJ�2��i�^�ij���}�V��R�JK��t����s�Ul(^�t��:��)�Þ���^$�����B����L7Z ��E�wOYZD�(�IX'�J��_�6�jX�;�Z���S]�.=� Ǽ|���_��$;��K깽Qt�Hp��t8HP���� �m� ;�A�F2�g���&!ߨ?�U>� TJ��$�F*v�3�'��Z]O%�A�t��o'�~{�lm�?'�/cʔ�Y���i�-���nŎe"��ѿ��9X�1HP��q�����@�%�ꍥ����I훀��F���#�ã���'�m`�H� ;G��������Ж���m���^�����r�C���WML�L��}^�M�?�Q�rZ�U/�b+t�d�X	�d��ࣺ�j�Zv/��H�-�s�Y�Z�U���=W¨[t(&��yz�m.�1�b8��|Y����8�y�L����n���sm�����`�+�x([s�|r�~A��?�#_�JӬ�Lt(�=Y�~�����Qd";�� ��~Z��h�.lV��[HΗ/WPb�e�7N��ESX���66�� �2�jcO��#�ד�����W��A��d�x:p/ ;v���Y��%NJ��|�ӝQ%y�M���}����q��w"��� ��Q�c�7.$�/ߔ�0VpJ���Wk�q���͎��A�����a�P�S��>�}�gm���Y_�\cB&�����o�>�P���<	.r�:�� ��_n�w�0�rr"��ON�?]�x�&�{8N	>���������4
&�TE�3���OʞV
(�X^&69C�MU�t�i=Ȣ���P���/�(5�����*&��g<S�?�m����8;ZM3Sx��/%�M��Þg����j:����%�w����(�=�BW��˪�/%c�['����[Ev�wS&�XO�ߢ�d�ç�v,�X�)��UL�����/�rj�Ro�=K">��ܡ�Zc��zLN~*dbM���$��G%{��|�r�s��q�A`�� jCK?C�U Q�����>�u0U(���
�nP1Eu���2
^\\sg����O��pX��t5�Q���(�M\�J4�����\UW��4<��j׺1]�Q�M�+rZJ��eMT�)A��� ��l�Q�Y��AN��A&��Q��gF��+߹s����A~�s\����b+ܿ:�~�c���R��_Lܢ���Ե��-��$\q�U��k���5��)���M^�n����S%3-K��	_#/��5|�KT���NO���::���Y(�/�?8�uP�x_&�d	O��/t�q�ݡ���LI��M��B�P�϶�t�d�~�(��2x@�K�hh��1��i�G�E�@^�o6�S�K���pB%z�Ӝ��A�_i���Xj�[(�ۨz�\��Ր���$:Gd�O�ؚ�����O�;���+�0;i�r�����$�vr������?���_^�ǭ�~Y�q�_]I����*��� �;���b:���~�H���i��������Q��X:uxY���mG1(�&�re]]� c�Z��vLV1�`���-K0�ݙk�;���@5��Y�#"��Q�T�P��>/�!ך�I��S/d�Wp4f�L�P?9ZA��5�߿Och��I2Ws'��}�ry�A�ز�\���^<`��]�|�����Ѐ���_��#��Qz�.�a�6	����Տo
o���iTO�n��(�ϣ1>X�W5��q�!��6x��R��|.5uuܵ�W��Z�E)��֗Է7�w6x��AP��of�,����ҿ�=�����T���3�lI������o`�!{ڦ�f��)NM���9H�B�u[fhuM�H��o����-�#��"4�^�,�9�=�q��".T�<'����F+e��dee�����F7,ѻF]UD�D>d�mOaʛ�i��� [�*K��س�j}�%�QT�M�� .�f>��Z�����_�(s���l�/�V��GZz\w�_oqB�^	��w[��0;%�j���#�"g�Y[������t���z����i�	�[������W�`	�f.C��kr���E1�7OԻ���5ʌ�R9�_��>'����L����42�C/��/���@y�ț���ܷy8�X�;Q��[8��`
L���j2|Fy�*�z�WO���D��-�5�qJ��-7g��b�S|�(���*���>��jp>��u}�&����A*���l

�@Ѧ�����/8+?Uݜ�l��,l��]O�v����R"G	����by������������@Q~S��6wy���?9i��Q�>_���D����K�Hd淌s��( �/_�<��NJ�a�3�--�Yf3��:l��%�5|p�����ᆃ0�+Eo�����w���k����8Qc�G�d���E��m�M�6�D
t٬��iG�eY��m^��T����l
����pc���wf�g��qH�����̒��oP*�{T#�m6�f�������ԗ��
��TF5�=��0����lbʢ��C^�y
��n���Y�-U�f�k���E��@��(!�����En^{%)�Ȧ/��=dny�k��j���6@&���묌m0��-aoq���p�Z9G�ꦦ��P���E�TD�Lo�@@��:voy�*�ư���eq߁k�ƚ�]8A��Ss�i_;ش�]Ա���`B) f��X��W:�#�us�Iw�����I�ɐ����V���>��K��'En�W��c���P�F݋� tb�_�H�2	ZwϠ��L���E�o,��¯?�5�\8oa���?)$���2	srr�E�A�v��s�R�׬�g���ֶI���F�R�sj^Φ������K�L������;�a~Ή��Dpپ��Z1��崟,��/�jS>>��Y+h��öe��
Q�ȜNg�Y��������bzL/z���t~��� ,y��<����ĺ�{�+��%R�� �?+�ߨ�Q���nz�9�M��R-�%=7��ܶ�	�F����]G�o� 1�4�vo�����U�����H�i�[�F�7�h�f]��LZO�Пdc�۝���vNM�y3o�2�+Â�N������w��0���Q7��Նa3�п�,��x5�Дd!^Q�>S�F�[w��_��ɶ�ϩ�7�P�l8IR�y���y�:�pr�DJ��UՏ^r��z,S�0tO���J}�lλ7��~��M�aıX�gyp�'�+��M���&m�[��@���B�g���'��"ϴw�j;�о(�X�[���v��k��8���l$n���|�ić�8�l��X��?<�rx[��@��=8=���C(0E�������ޭ�1�\P�?:h���zἺZn��*wn���0[���?pJě�Z�v ���7����d֏8�;쫙e�ȏ�����*暎̋/�AY�� �u˛��q��`|����L.i��X��x���ʹ���A���p��C� ��߾!@�<�i��:'d:A��݇kY2����E���n�V��Ug�|��j^�����?��������|�����ȝ7����_C��ӕ�>��ϑ]KZ���~�&t �wX�7���ɯg@����f
�O���!Dn�nU��B���A �в�8�!����z 8��;��<f&�}�J�L>�F�Gp�C^j��R�B��F/�]��C�%G�rvL���^�u�f���W��+g �{R �T��=��J$+�O ������	�b3 ߜ�h�~m�R�k�f�Y�Z0W�.�f�=�(�\��ax}aa��>=��Z�}Ҿ98�^3�*n!3�i8�Dd����n�Uꁰ늁I�MW��F�xCZ�����}ǽkղ�lT�������\�3�v:W���� �����F��R1��#m`�P�<{hQ�"��F�]���Rb걺
 ��� ʶ �mj��� d�/��]�΂��8�	��=P�0  c����g`s@0} [�A_�`�����s�I$@.�Y��'����1Dk�AF"Ѡgi��\�p4ٵ����A��Iָ�&�a�7��5L�(����E��R�����8��K
���X�bF�0�y_��(���}#��0O}��0z����F�H����W�#���/���d�	� ���}ŉ�}�B���g5� F���N� r>�5pF�ʋgkMB��z�t8�8R���҅��z��#~&($c�뱘;Z-�V�ɠ6σ}C[Fwy�N�Z����g��ρ�{��F��,Ɲkmu�Kbm���$����yP�� $����/Md�E�wI�h�x'
�O�D���Sm��TL��^��Ec$]1�u�(�v��SvZ��ݸ�����?o�C<p:7��>��Pؿ�ޱ��V�=B"_�3�D\����	N^�ܤ��s���5�,ʁ�o¯�K��
�qJ�;-Mb�#I�y�|<��ր�@���Z�A������_�574 �|%	 ��;��U3x��f��2�㚭�c����v��2.�[n��#Jq����9�����\��[ogg����u��-W�-f��&#��r�D�\Ҫ������� "}wEw;��UP-�<kY�{��G�`��+6O�^M�Fҫ�e�Hw~�ܥ>Ǎ��º2cP��Y�%��Y~sp��ΫF�J#�(�ɥ�&�ƃ���q�O�l>�Du�|n�E��P�]8���e�� �(J���ݣy���f|�}��.��}��C�i�W�^'��@�b�'��K8�����|�gG����L&_���dѾ#�s��IVz)��C��|s�]�����R-A�|���&`f%���={�I�Z?YOC��m5���1A�,^��k�J�d��<��S����~�B��L≿0٭}k�3��L`��4��#����TDP�@����bj�'��@��kv+��h|o'��߸�P8E��.־f�t�M�]�����>�/�>S���g��/
^��ȫ.�&$�׳����75�M����bf����������,L�,��߯y�/¬A�(y�Q1�#���lj�b+\��|��߫F>�tΜ�A�WA�6Lv�Q�	9�O�,�jh������R��f�n��<7��x���j֬�Id7�/�L���p���w8_ ��r�
����f!��Kt.P��T������DANM�� �����K���*Z�޽����N>j*����\]�V ��*���p в��0�aB��xQ�_�x%�l�l�AT��uV> ����ߥ��Y*eRɏ�w�O���r�)Ȳ �..Q���3���7���+��GgL
x�������� O�7�Y�f�,M�;~7�jf�@/<+��mh/XN -���J~w&k+��/����Y�L ��pL�кش���qw����S3�V!p(н�
�q��?k���|����dbg7V~5)~��=��|�|�܍��?`���f{�K:�J�~� �*s��?�b
�BfzVw?Vp��2�6Lຘܖy6�y̋t�Zٍ���@���>���i���b7�ܜ/h�co�e1y��^��S�A(8�ŹG9�B*~]S� F�����3���r�SF�'�lM�i9G�!Ci�B�҅>A3��Ϭ�wA�.\-�_��Ȗk�h�Aa��S��l�2������~"Y���8^�<Y�2c�h���P!��"�@Q���B�w��Q�T�ư�$σ��y������ܮ�U��ٌ���4����j�d���=H���A0w��%�Y�p���6��{޿j�� ��]E�&�LM��d�ʁ�s�u���{ۅ��b1\t0ϩD�<��㨙����ځ݄�$ɳ
T��V���/vE�t�B�~Cżw�$ll/���B�	�7�9ՈIt�i PX .�y�}nOŠ���D���-\���+Z{�ps�.�5`�\��*�S�נ��Q��0��D �g�"��뱒���Z�*��;��V��8��!q] WW�U���_��A��Q�|,$���.qn���M�ۄ���Fv�������f�ފs�:�!�X~&�|7����x��ƿ���Ӌe�<�L��K�G�=�����ƞt~R��I��F�j����UIKge��f�=���uD
�ޕ���!;s��ȅ��ѠW�����Ye�ʅ1w�	��+�� \��5�[�� r�5�#?]��?�@o^�pS(���z1�A߈�����"��*�V59���˾ɞq6A�?��ȀN��}/����)38;m��"�/���u�	1��@Ԍr�Ŀ?��"��lhg��hm����8<LGuKo�N�s��'ͦX3I��l�O��Civ�@9$�6���@���Pp�K����?w�9Ժ�Z<@Honm�>�ꕵ���աC��t�+n�t���tm����Yib"}� �pV�������;��)V��C�Woݺ=2lKF�P�m�I4�S-���ܛ}^�}�amaN����D��JE�����z����� �m��Hqp�ߤ}�u���-3��Z��| �YD"ߴ���)5r!����u:_2��N�9h�3��=�V��M��	�x��"�S���AeWL�ő�8�MInáȻT�va�v�R�J��@���(E3&���LζB��⾏�l�,�����%ȍDƖ�$��p�8~��QJ4BJ����3���Ъos`��n���Ň2@d�-A�9����ç߂�Q1E��%*~�|�ϟy��ʥS�'t��8�^�+.�d���q%˨۩�� ���r�*k�&ӌ1[C/˛�g�B���i�R�T�* ��j>������6&�v�ڳ��{ZS%H.û��v�r/���h���S���/#�\��Df��^�t�ףC���9	��>�d���싒�>|0M*8���{�R�4�Zrs'��y�p��LN=�yHi�N��bֹ��f �t�}�s���iHC���L�R�w��p���&
�����足���y��/VWr��oU2��χ/��Q�4uL�o�������vy0�~G/���!�����VcS÷0����֐-KH�1CW��7�$4!xR�*�\I��DK�wH��B�IZ��g�>�*�3��޵_k��Xg\�qa򣇚@P�iH�K�ۍ�/��!�J��_fo�z���H�a�y�����w���L+cRi�W2Yu)��}���¨� Y�gV�S�=姗���KSݏ�߾�=[��bm��k��<d�R�d�E"1(�Ї~�u�$ݹmC3N�=�L�y�{�TӲzN��c����*��W�n���f�)k��J�Z\��P�u�Yg-q�����V�,����8I��������ö�[�>������jO=Ş�,=��
i$ku���O�)�W�iǉ&zeg�1d�|H�N���PX��<t<��ٝ�_�)���7.�4������F���ocF}t�:K2Є���4�4�j�VZ6�Az�
���M/���������R���*��d
MS�=:�Kk#N�pVl�T����;��Z&���?~@9�x^�"_)�AC[r���0E��L6��!�ߓ3�`�YSb�H~d��M��'aT����f� ^�����m1[9�ǂ<k���$�5Bއ*��o{.����Y�:�1=��o���}��3�'/$�]U6j�E{�
_�|~]�xs�E�GW�ַ���^;�^;b�>�FX~�S���s��DC�u�U��� ���������ay�D�~�x����mcէ&�ͫd��W��O.��\�>��+?&�/,a�������A��c%&��>^�E�����S�Ny�d�4�2���	W$�x��ّ�P��9��Z7�?x�jȺ�mE�2�����塋����������G��Z�\
=�R��U4f�Cm�o���z5����yHQ2�:!(�v@Q;�|0�_|����!�;*M�-��(�-��C!����H:P$��Ӭ�?���.����
]��7��V��V>7�[�(�}+#�3s��%�}$r��$x4&�uuಊ�z�b�N'H�~��iz&��d� ��S .��utsd-�'*�uU��ˎ7�\��e��l>kY�C(�ds���yW� ]I�}�y�acH�ԋ��8N�Kv!5k����!.�2�.����=��¢�[��4��]W�@���
~AG�
Ɍ�"ъu�܄���ٚt��%-Ä!�!�&�G��˦0;BL1�FE(��B�}Z�C������;3�.�)$�Q7�)��6�]���V�uy�9�B��aT�<4[��������L�n�]��(��;�w�����혳����xڑD��p�������ֆav�B%�"u�3�G��CN��S��%L��c��%�hh���᩟�y��A�6�����{�.|n�^���gD_ن�2�"���=jH��ԋV��{�x�yQ��w���q��C�Iw^�B�I����Z�X��Ʉ�/�,x�%٧B�)���Ǻ:���7�y�N��C%�(��u�=��Ph�vt�;4f��\�f�S�A�y�������%����Ȱ��I�S��s`7���~t�ǭv���e$9�����U��= ̟���������B!�7�Q%.����W�4�u'|>7��=Fzl�N����N`������B���	���/_�jZ��=dۊ�1f�5�Ǎgn^U��>����
zб�]��g���<�� 臇��n�>��	�hfZ�уҼB��i+��j�7�����U����<��	����^PZK����� �;鋯�։Q��7S/*��B|�}RΪK��٭�2��Rz:ZwH-%8�\��3�Ҳ|���?���%�� ��ͦm��VƶM����������)��PH� �MO������ۼ��ǉ֞*�ރ?�n� +[�N�i^Y�H��ܐB�����~1Hꨜ;�<���F2�c�z;S��ǍV 9/3����X|:J��聙�93Ҋ�:�;dp��y��DgagW�w���x���*'X��F}�۰5�<^��|�2��mm�v K���{�,3������穜?bQ^�i��¹�����kU��N��$�����V�=��I���3���Bx�n��R�y��P�ҍ�'�i^�*��ă=�����eF�Z�N3C8XFO�hXY�s">�5ơs�Љ�<k����)�c���y�f����$�D���3Չh2͓��~��N>C��YA=
*��{�A�Ba���k͎��mAS��M�0bY��L\���
TXMK�YC@Da�v����y� u{��eׅmN$J@ �cײ�����/L0�[P�d����ᅅ����Y�%��S�i�k���S�� �*����wH����g^��f���m^���y<^<�-ɬ�lԟ��gB����,7�{�3,��64�@�:�+?���H,�E��%���B~ ���^��\Q��̉��Ϝ�2o8�Y����E(Q�X}M�p-�b�����ؑt�Ot�<`�,��������fW?Iy�#�Ĕ�w�6*/��xT�!�Oo������P�j�˛�w3�!�g������n�ߙr��-Vݱ�7��,��u��Tx����0-1���`l��\y9�O0$���[��	u��"{�d H*����Vr����3�q�a��)�[�O��_14�>n��%c�D��%*��Z���Ԗ��0a�a�BF:0���]����E9�8���y���'��a��P�d��'��Mƫ��=:��(���m�55�`�ږl0[�͎%�
b�0��y��Sv���@��D;6�f�g�n+��Q�η�X:�1�����k����v ��!![�G���]0 e������N����B�4�Bv<z���DH�LR���u�g�B�����_���3�<���=v���uJ0�"|'5�%�6��ZȦ|]3�����%\Z/��F�eg����>�q��D�à3����S��ۢ^PK&�'����Vח���t�'I���'r���j�zk#��Л �������s�X�<?� �c?ƣ$��m�b�;	��e4���ۼ�a���k��[��=r�D��4�/�WL �.� ������` �Ѩ��䟭}�W���)�"N�Er�,p��d2y%�Z��r�n���d��(�3�O��;��:��!|�A��k��Q͎�-7Gd�u��g�!���;M�+x�1�~Ƃَ���r=xBq���_E��Zd���x`�Jؠ�������eᎩ�si:�A�u�=�����t�Ӑd��=-Z��}�q�'��m_	�8QO
�gbG$�ӾG�P��(�	^"�����v��,�r3u_�ǿ?������I~��=P�2�
~[+9�b瞞�`�<"}�So���>�T�>�#���L=�Y;��/T"����cN�W0��A���!`�v���nJb��v|9�;�J���3�..r�Z�ր8���uÈh8|:F�[��(zj��|�'��#�설B���B�N�7�.�8.�V�@lo��b�T��H���i?ğ>�ހ���}zm�Y2B�oC�&�Tr��3
��Ժ:�艃��G@�b��A�c}�܇N��d����@��(��f��ŶՔ�#9������[���An�&��Ծּ�f�w�A!|�����z�0˛F6��R���e���v�1e7��q��Ϋ�P�O����>l�$�^���ӵI��>{���g��W�)~*Ѭ 6�m�
�퓋� L<C�	ؓ�o���<eC�><=�r��yC�Q&r����߹Z�h���n�ޘВ�3�
�f�
�L�kf��/��4$�-	i�?�d�n��?������zXA���B�l��[v����x���'IĖ'k"И�y��|y���(��٨SE�����q����K�!���P�
͞���[��2G�s�,}�*��)�&!p$Șd�j�;����lI�4L��{�7���lѵ�8�蚛�}�|PŘ�{��&�>��۲�����
�#R^����0t��N�w��:��.3o�ՠ��`�� sP��d��6�d���5$�'/
�+Iy���+��Q��9 J���b_���o8a7�t�ȇy9_�,%�.��	2&��R �WDfxȬ��ɓ7OK��1I�-db@n]y�7��B��p�<tz�"�E.���1�^��]�k�t����Յ虎gY G�tnJ�o��"������i�� `e˹l���da�\,[��+��t�t.��(�7����(2����>͆�����Q�C�<�a��е(�e����K���-ےxǠ���45��PA�ץi�o�� �����|�ĠR]X�&e06��{Vo }���#�-�t�	J?�*��&W������TI�����w���=`�(���Hs�e�5����=�O���e��&P�py�	[k��G�M�V�L῭���e~�GA���?�ªk���u������s6K8�r�R� �q��]� zJ����yK��[��<r�4�h�t�9�N�3��T�&�Rr�+��PO������ ^��5/�r����6t�`��U��Y�#�`�Z���Z�����l�2*�l
�=�)P?��8M[���)P�da�����x?O��O �������Kx?�c���V¹oa�@]���Qo��g�婋��N��S\�~c|AL�����|��5r�f�A/"�|I>-<E�z^Fj��.|�ˉ3�-7���O��=���O7&��������lA��¡Y����?
H���n�./���[C\O�FX <��Y�z녭��T�wå��.S�Rr����4x�E��Ԗ��W�]�6kf<iƿ|W����ᢅ�?�߆l�M�0{��Tޅ�Dh��~%��h�k��Y*��PB�"���I5i
Ɏ7�_qS|6]/<��g�h��oڧ��28��������N�����#�Ջ��Y�&A4fx�a���>*�"�(M�^"�.}r�jb��7�)�Ky�d�0�bz���p��j������p^��MH7K�^�J?�B�9�BJ�D�E ��X��\kk�π�d��z�$��!�g4t[^]j��a�|R�����t_/J'������b��ӕW��ҧ~4��{�>�Z�dѝf~t�3F�I�6Ki����|@ ���z�����9�N���jO�����Olw�

�t�Iֳ*�G�X)��gDq��K�<�,3T7�[pe�0�}��+)En���C(��ND1�l�!s�2՝�.�e2�R���:+㣨�!����d��U>HW�@���1�z�KYӾ��=����V5��1M*�1��s�y��ֵ޷���۝ipz=���!;MC�,��_��+}hul��c���̻5K�����[���l�`�Qs���7g�hy�8�O��-l���~@�y�=4�k|��f���}���F!?`�+��h߁�Z%:;r����d�DY��v�q���������&�ǻ��<BI��IBc��B L>�U�>_�sbs�̊	(ϻ��j_�/7;d�l�����U$�
�܊s�Ƽ���aڝ�-�a��!�P��R����z֊X^�}Ⲗ���W����:1��a�K�9(�	<�^��~�5fR���E>�F�`jHlK}�����0i3�/NIx�&�-#��
,�:��\F��?�\�~�xl��2&��ݳ��O�Ig�a� B�p߇J��g�_	@���d��V'Fa �n$����"瞚���s��F}3տ���ĖKV�d����� �
Z�E�m�(hN�^(:�X�����k�(���i��2�X(Lc�9�A�@*�57���_�(�3�3׃�X�;TK����=oU�C�C9��'_J�����b
1gC _��脙O����9� �i������dSP�9緜?��Q�0����!���B���}�n���q�9�R�m%f��Ӆ�΢~�M�-j�a�Ѯ%�7�c'L�a�#����U�2dih�X�������f]���E��oxf��1�Yg���Y��o+'���_�@����eq�P&���1^��t���,�"~�'y�@���/'[c�UL�L���U�7B(׸$= ��x��݊;P����`�?�[X���]�'��}jV|�M���}����e�Z��}$�=GP�w���L�����t&֡}���L���{}��l�c�r�xi��gf��nH"w�qɝ��|S���s<&o'ڪ�Jj��S;��nÇQLyM�*k�""0�$HR��r�1O��lOՂ�-�2^��:�E�St�=��;���%Doo����{���k�^������l����;�
���*ʜ�������>�gDF���j9f�oT��,��7s��9�@��~�;�ef�(�	���j�F��X��|�dҨn!�@���%���դ�����E�K�� 4X
.��d-�k# �S,va�E����6� ��iVZ�	,�	}z˝��������x[qB�I_ɶ��}I+9'�9y?������О*���+:q��X��"�l�@�J.� �v~ �Q�}��:nǹ�_��j4y7��\4��o�7���9* Y�$LyGuG`�M��򚆗��iYp�yUc���lJ6Cx�(z���}._bkz皮���ɏLG�=�p#�_��Y����r����Vl|1$O2�I>F���5�b����OK������R���-M��;���4}ӕ������-��5����?��u+�}ezB�zU�"����5AK\�\L�ઃ���įlWh��u��Έ�<�U�k�w������8Z7��J�.�2�;��]���;��<��e�ʹ��D�<� YPw�`��o��z�`r��|+C��N�R^|�͸���t�P�Z×o+�$Us�G�{��f�s�����7t&�ѤkĳC�dOT A\Y��lMlA���*ڬ!��[*i�q�v�;p�Çz�W�3A�9/5Ch5\C��ً�ժ�AWn���^9����\����l�5}oxT2칶jOa��-�",S��?��n��3s��~�K��z��@��Y/��^��z,s0&���}%�}I��W3��t�l��d�h-�����l8j�`�TL����Cb\����u4r� g�ު����/ G?��m��ŗ*>Z�p�9�>/�ޠG6�9ǡ�"�F�1����/"��cp<�{b�E�}G��0\V�X�=��'+dZ�h��.<�z��N��g����h\��G>�lM���F��*��:�S�W��#n��As��	צ�N�Ĕ!G(�9O���N'���B����y�Qy���|�'�7���П��Y��~Wt-F�\�����x��s��ނ X��B��I߱�i΍[o���W,��/J����廖d��s�ĺkf��)9P*����r���%Bȩ����"�1�L4��?e��$s�|`s`O�L�WΫ_+���鋍3���$'9�KI]�$?7�(�t�S��-��EBc6qnyZ�e��9�.wv�ϛ�h�p;�Dv��l�Ls�Gx?����Ċ�j�'#�I��nw��l���=_�x�gn�~C#CC���1� �d�R��>S�^��4z F�i�Y`G�R�y6���βyXY��n.P?/�d�f�u�Ċ�59
!V^WTT\�)������%'҉;��bxs@���Wֶ:j���Ї�.��
RKTkz�>�G����Ƴ=��8a������&�'�Bgo��2;�R�*Q�k�wU�9�bj��h�o�T���~�H�6{��H}Yy���^n����.i�T��/7O[8���;O Y_	d˥|<�f ��w6,a撹�J�q�@��9��P6�4[*ER�q` ����IyQ���
��Ԃ.�3��<\q�e����^�1��xBP�d���s?zP���-S��D؍������<�x�iqJ�(������Ym���l|ߪ?5鿧u���L��KT�IS-��?ƍ�BqU�F�x=x{�ã���t؝,�|FlNz屔?�'$�U['dcy�R���N-i0�\�����j�PE���T�b4�X�@ٙ�
,v�;<�j(�g���?�qQ�z��;B"x�\"���*��߰)-h��V*�çXڬ9�l��Xn���~|�f����iN��3�\��7�b��h16}�s.�у�s�z�֕�e2Ag{aǟj 䎅�#7�U���s9�F���Cq�"��ǚ�l�<�̠�d�b�W@�e��g|�-p�!m0��jMC���0?��Y�AW��������I	���Y"�t�FҦ�e�������9���.\��:�
|�+ t�M�ɦ��E�̼T���Zd֒�j�`�ӷ��Z�m?�������ZF&�M��HގZ��!�P�g��5-�bw_�*��٤���O*\�S�J�.�D���qQ,�Ċk��(��\����G��ګ_q[;����U�P��iBO���\���D�Yo�;�t���~Q�5�Am�S�����J=j-��:�Lq�(L@�5u��L�p�Qܘ)�=�����	��Rh_#A�7T�ò_�~�|�gUڼ%K�o}딬`~�z��>�(�#g&��Y��@�T��9ڎw��5�l���2����Y�ө����z�#
ßs=�x^-ᤲ���B��W��F*9�µ��_k�{I�@�gd��Sx䏀��WM�
-�5aw?w���|Tآ$D���ǧ�5��~�����'��@;
���W�0�q'qKP̳��[m��(���өT��FN)s���C\{4��Pe��$P�������b��H[�WE���
s�UP�������9Ǧ��cū��&k�a� a��˗����%�	ưm���|J_�J�-L5�SQj���+���AQ�m�i(�qCU$���V�et���hy�����ń�#����ac�������</��I��7���S~I4Fm�E�U�r��UDHWr/5Xդ,iu5�AOL_�R��q�nD�����Kr�����C�[�E�}��C�� #����-��2(�))���A�F���i)閖~�|�Ϗ�������^k��u���9�W3=b��@S~�6r+�B�����$?J�.��;U6^a�jǽ� �����¹��ZZZ,c�f�	o*.�c�_�G���ºɔ�>�$E��ajG�֯�z-I�:�0G�ȈLV����)٢>�<a�%��T�Pg����ఠ��qܪ��m��c��xPN��\���:�h�����]ԲiEw��"q�������0����!Xat��j�G%�T,��~K�=&�~�F���%�5J�'�h�J�fHw�ۡ��~� ��L%��$G�?�fk���$䁱���{@�f�.���ǅ�O��FF�����3X��Y�TTx�>z��G���}_dÞ��)ۼ�����Xh`X��o�JT�gj�������"xܽ�]���9᧡���o.��n�|��{��R2���}�R�������-,�0�5�٠��_o�0/�T�t�)�¹��H���Ĕ�r
r��4�R�K���h!�~����@d4�wvv�G��&�޸�t`©���$5��bU��j��Y̶�(;������׹�=W���U���m("�6�t�ѵ�4I�.�;E�\HgN��m?��*�� d���q�[�W]����B����D�"b6f*p��Bc0�ƮL'l?W��6���DB-W+�Qn.=���r�D�G�rq��QVWd!�b��8ͼ��|8�!�۷�����x\6�Y,�+����w�`ܔH���YkVjrr�A�f����17|�+�gҢ*,��SR~��!Y�a��y7<�����?��l~��2��U1y�M���H�3�c��f�g�D���i��`��Z�lTQa����o�;�T�V�D~.��S�%��iog{[�#��A̔ �{
"��e���In��i����kt���1��/�2ĊJJn����]	`���C)�oNw�h^ki�bx�f���ҹ��*ϘXo1�We5o�s��s�B���2n��lRҠ���+��լ�͛dE%�k����Y�X~*#d�KJ�ܻ�!~-�RRRi����<LQǱl���gKyT7V|�7�a������MsS&S�М�܍�A?0�Ē�QW���5�k&�u����3$$$���
���(3�}�'�Y���S�Ǵ;$p���
y��߲1���WU%�q�����_]_������'ZJm(����񋘣�`P��9[B�~���M#
�f��Z��<f�֋E���GN$���S���8��2��PG�)-ݳX �+��dT��{���8�Xk!]Y�vI���/��[,�D�e#HB���z�͉`M�$�ð�H=ruEIp\#ll�8�f�Ғ���R(L��#^�K	����;��O1_��)3@������*#�Vj�pG�@׵�h�^�芓�3�*�L�+)y�դ����cD����D�Z�b�ϫ7c�,QO��Y瓰��b��c�xUx��mt��O6��˯U�{������`H���<?=?G0>T��tl��1H�A���B�w��.@��}�����N������fL9��F��������AEtIIT��4�4:�Z�vx��@������f�C�2V7$����W����2��Cڗ�����^D=��b���+��� ���D_4�Ћ>1���"�C3�i��+��o_�ǟ���ӭ+zMR����=��K	�f���m������������/_�\vJZT焇~���������H���^A1�ܾU��x�'���kɺw<6�sY�jڥ�L�lzEp��Fs�0�%?rDn�"�6|����$V��Gf�����i�3��"�s䙘%��A���?yn.�V�:J$C�Ss������Ї�G;U~�v"66V��ּE;D��b�#H�d��{*	_Ja�o:�\��Wswf�P�nn�����<S�jV�����5g���׬��Z�u��	B��O� ���0?p�
�1xyy�EM����IO��DQF�ujKh�b.�^��K�4���ᮡ����T�}Et@���v�n��y��|���Ъ��2���F���oѣy�mɞ<ל�9��e!��ΐ`hh8��@��Ǳ��t	,i�5��:������w�o( �q�4��=�l����G~:�E<A[��SfM��mo���c�2]�<iH*�0d�r,(��&��AJ͟������#jmc#x�2�b�O�FZ�5���ϨGF@y��ʱG��pA޲�X���M�$fR����&{����sn�8�f�IpS����N�43'�;e2211m;oCȻW��σKJ�89���҉��IJ��2	(}0���ι*��x�b���g��G�ɚ���@�U��9��q�T�Vt�V��J��e^�uE6g��D��������y�=I�t1gPHԜZ�f�M����N�x�cY���sȼ�WdD!q�v~�e�"g=0�����O�~_{c���Dq[�����1j��5}O��n�Ն�"�e|�X�Ʉ���I���L��j�.�:��J��%V�`A@�N#%fT8Y��:Њt8'� 9iA��[��3,���TP*�R�/2\�e�)�8�%�n�(L��M�[O/���J���&����H�ÒQ��}���ϟ�ݱ�F
�q*�͗�󙉅3�;^~?k��\$��;�3z�]�A]Y���J#$�V�<��`�ZF����G�m�`n*-�.��͔��6?=�M�Ud���h��.xQ`�$�Љ�z��d����"� C���_�=>�kt��K�E4"vzz*�Ljj	�_}@�����f�*��TS�H���b��U�p6���P~
?i����� �s7&{���yqZ^^���E��/���-��m��@sJ$�i��`D���৓v��&��]�?����HI���s**����\(Lf��c���ܞ�� Y�aw���8��qw�G�Ak��B������_J�GG�j���n�G�5HQ/�Ω��a��'�-]��%��H�50�[�[��.6��r`��0"ĳm1y�\�.߇M�1\w����D��v����tQyv󢉌����ZE�|�h��}��G5hH�M�,K[��P�]b�-R�E���ڰ��v�3�^�Єܶ)����x�Ù�]����ȞF��O)��?8p m�h�F�e��{�P�Y��j�|�(��EK`�	��蠄N�]r�P�;d�e���OY`�VӟQ�����O����\��4m�L5Q��C�/?���u�e-N�˓�:l�X'3y��}����E��b)�����}�%.L�t�m�Zq���_��Q�|_��>t�*�@���O�e����)��5��O �Ȇ)���[7(��'�'��6o�>�rB-޿��I�R9c5��D�4�V��6~V�|$��$[�9r�
M��d{w7@�,R��)����z�!2���\�$M&ز��"�I�A���W�P����)-.�	��x5w��i;˾�\R"����[�����jsy����JPMI	��2�x��ѵ���H�+��g�[\�|��N�s�� �_J�А�ʛ�SB�0"�ƿ�%ł2��F�l�����>��w�F�g�%�1m��gO`��a��O?bS���8}�)�b�����+����Y��
���3?ŘQ}�Z�]/z�f~H!��;azc�%t��o�8��X�F���R�y_"�c���7CLq�Z���NRv��""����tp|3)z�D�iMo:7�GWl?�y�BgJ�����|��ͱ�9��
����c��D�a�b�?�������n0�=g3�y����%:R�eo�
�^���n�K�	/�ȉg�t4��$�n�m$05J�����m	bcx�w�H�T��?�V ��BKd�,U����t����k��!�v�(��`�1��]mc��Ӥ��~�l����Uhk0%is�}��
��l��i��Ą������f��weUՑ*��X@�@���[Z3|���W����Hd��/`�ߝ3l)Cs��b��eX��㸕���\Rr����a�OVNn�L��%U����S΀Ĕ�kjjZ~�D��՟�b)N8�и�Yj,��u��̊�D�w�Kdt~�W�W�3�̠�jVa*�Ԯ��NT�h��҅i�W�ag5߾�|oBN�Ѫ�R��W�i����W�Hs~��G��o'�M[���禩��*9�Ƃj����	��̈́<������K�[��
`U��?6O$K
[0._\綴P.|,��7ŧB7s��t1Ml}�*ݚ��g7{S|��$��V��)���mf>��N��"��O�~[�����GY��)`W�褬�;���z��-O�@t�I����.�������Ց��4언��@*��e
���R���V��l�D��NP����
���Eb����-�x/��jO0S�d����˸��ș���-�_"#$�Cπ�E����Sŭ�W��
�\5B�Y)bw(y,6r�����k��fnL�@�Ј�47�=Q���~Mڵ��jt�o��EP9���%��#��߽���Ѷ-�$�Ÿ�	�f5�(��8Ŋ%���j_ϧU�>{��I��*�
�5�l(�X=6#��%�0+Pj]pؔ�`��wXS�u��7��U/8x����Ii���K��U��M|� ���i�����~?Zv:h0~ӫ��l�@���C�n�5��ޚ?���U��f3��rvмH���Q����`�#��� �cQK}��'
�.}�y%$&Z�������Vy�w��k&TJ�UI�� �Ѩ�� U+� ����
�!ۡT�}}h 0����q��{7�����޷i)��$2�c)WWW�<̈́��T=v�[�����#�G��RTIe>�>)���CBz���mD_<�q��O<99)��|7h�G��}V�����;����� 27����v^0Ȏ�S��0U��Ib������ĝ��UA���6P,�T�VCO'A*���y�ЄxQ�x��d,t���))��:[�?�'c�2�:U�?5�MIA�_��%��2�Q�h,_�ߋ�-�����L�{�f�{E7*!r��̑u��v���O0X����νʾÇsM.�O�6_SDzf1����IH��7|��|�
�Ft�R�UA����K������qW��I-�aH�U0�G�{�m���wo�d׹���Ԯ�9��\�ǲ��(����`A.�YǱ�C��&�{����rq�^�ɚ3uo�O�Ϊ^�7���TS�{��*���#���ػS���TX~�=�ġs�9r���TMW���ٙ��Z�ڜ�F��+���������;O�7�9�%��	��qZ��q��8^����"����>�����X>�	�Z]R{M�Z��2�M.�h�].j�s��2W�:3f���t4��ڊ*�(�Jլ]ݴQ�_�X� ��RH�����b�/��G�0(�r��r�Ѳi.���Q��^��
>%A�B`?�,k!'����y'�����A;;;n��&X)EJ��w�\�b�e���P'# "ڭ�qi���cj�~�Z��a'���p]as�,{�E'%�H9��d��X�T��?`�Y~@�{tx�Ʋ.gVu���|������wE��C�Sl�C��FB93.^ �[��O=hu�t�ȳOcu9�U�G��Kfqh}~���z��
�o�aaa6m�?����C�1�q��$���wd��UT�XN]G�q����//��o�@�^t�I�lF�+n�(f>�3qݦ�z�74d���f�LRF���	v�/>c�o�0/	-��!!nd��ǃd|I����󑥀��3i�:srJU��iʒ8�)Q6ś�?��XY�5V$�e}�
h�#��*�8>��[���%L�u�5He6�W���~�KXXXhd�X��;JYY�=}�s�kd�A�y�أ�������i�wn��gI�1�:)
��4�m�0�?Ez�R������Ɯp�ǲ��E�h�#+���J\8�<q�����:3��y;_3YrS�Z��C�:��P��}�&���^Л���l�8͒�0
��t~�4��!�2�u�&�樵nJ�м�'�J��5.���^������Z��������������p�e�X,��
J�����:8���'#�`k*Rlsm�"A|�c����-�Vz�8��#Z��x�����}O��Ϟ������/���Z<=������'��U7�\�����֚/7�.//�)�zOD�V�)s

~|>.��GF&�����ԕZ;�������=9t9I��z���*�~����5/nHHO�������]G�0PsII�]Gss3�."r�uك���E�ժ��`B�[���`yצ�U��\�vQ�b�ذ�J!+L~�D�<>~g%%Rju(:8hY�a} Uءe�>#*
׹���p*�Ŷ�}��c�m'K�P�r�:S{�	���~�w����;����q^e-;��"	̜�<=����l�d~ۋ�4*�<����±�+@X?�☿p՘г˸���ݭ�)b���z>K�G�^�g�knk��8;:����+ P�v�����U�,�u�X,-��������N�"n�(�r��I^���iW����|��5)�x�>�%2G١^n�T)�7)c�}������\��}���Sd
�λ���Fl���v*�I�������o��ڨ54h!	8J'e��_���f�IA*/f�U�,����N�Y����c%us�h _QP�ˋ��W�s��-����å�Db�|�r/>��l�E9Cԇl�s���Oԋ���<�Qy� �_n�[��n������t�K�����[]=��i�C���F��� ����y��iii�1�]Q�9L6?����OL'����y��f�o��"�K�վD��̭�(�b����˼�/�U�%Z�	,R��"�b\���ʼ�TF������ ������=��X�!��М�C��ҕ��e����?\@M���</�Ɉd�a�����ѱ�ktZ1��A���ɨ�����+Wż��=K@�d࣯P'���Z+J����ֿaL<�!t2��r��)��ȟ�ru7�;���*�C.W��2����H���O*��P7g���އ�X�<kk������}Q�ʽ��(�Y�#$r]��8���JW'��n�,��\�Ʋ�a��1ChG�T�f�,K�\h�ϟ?W���߂U/��)���{��`��	���I�w�{���h����D��8��=�z�:-M=OC]����+pe4��>������dnnf捍+54V&��݂�tU��GQ�ӡË���̀�~F� 1_!��_���A49ǔ��!�{̐��БM�~�y,�!9��d��H�0���Dݹ�w׿����7g]�����i�����p��nllH"�	Cf�=���iE���H�H0'�R�ƾ��Oy�b����Ƭ�X^�L+M��;IIu=��e
�/��E�?,v�W�tb˦yLg�2JR9�"=z���3���Yg0V��bU��C"��(�id�k��pQJew#%'�ۦ����k9F��}Ş�7gb��<R�p���߭���b�~���x�ͧΚ���2�����
����ʾ�}ο���T�,�z��O��d���7��y��`z�!V^Qad��U���y��ߞb������Y�((�o���ų'���H�j��[[���ަ���x��jͭ����G� �[���ot�e7��/=�w�y
�w����5�[+Ds�za�S0!�-!������oooŇ��~*���b�k6�4�f��G�/80WT叉>rr$�(R��taa�l��*yZ�t�P��� ���$ث"���|>5�pn�:cm��1���_JJڟ��p�>�g�i����|�j�����H4���ݰ˓�yˡ���v��ӉO��#'{Ijbcl"z6��<�"Pw��!�j:.�㇡0���|��Gq�M{���&W���7˯*C��ͮ.�Ac����f�@:h�
|\2^�Uq[O�D&yߞn���i�+{rN�����%�� -$RRR����B���c�ʊ	��Knmm2P`�T��Lb��KJJ������+�}�vk����<@��L�Ϲ]SN��������H���/_X��믺�el۝��os3G��6�7S5��Ҳ4222m�0Z��O���k���8�G�P��͠�KO'�˖��8�XM��'Y��:4$hR�s%�Q��h(L��:��Nƕ��Y{at��ʳ� ���vo߆ ��>^���D��eC�>�	��;/�&*�$&5YBj!RLt��p�8:����w`N?���߲��P����������|����ͽ�h��%č��9�)|1���O�J�F�NW�B�O�[{>q�4��Qſ��hq�|��U�
�?�����oMϘ�,%X,�zD�FG+n����,�:�����[;8��5!�ș+"*q*��=nm}}��h3|s22�7t�o*;�Q�֗�榩_B�>��
��'���f�܅�X�B�i�Ĉ��3Lhn��		�\[��iz������5�V�(�r�FБ��֮�u����yi��$�9����"� K[����gm�?���p��xv�x�����4@�J`�)8�ssx���w��ȇ̩/��~ͥ�A1���b�d���W��-�/ ���e?}(�/3l�����SQ����).f*�gcg�B;pz��.X n�)����yYY�
�踫��Ơ�@��
^(&]h��<c�gr�e�!~j���PSC�s$KTox`�d5�w)p�ɐg�xq�D��������*��\1��q&8�����Y�9��f�����/&�ʅj�J�xӉ������|�枹M�]�.�D��%_���5�����?cW��߂q|[R���MgSz�@ō��X|����tP��Ui}=��B����2�5v�G��@'֕��;�?Gh{F�H�������[��$R���q2� E5(AϿ��z�<��" �o	#V��Y��G'�����mlm��.tӇ,��K��[�V���>	��:��g@��ƥ��\2�ZK���5_���,�?��^k��*ϓ�!��<�����5j+×Y�0��Σ՞ܢ�p6�Fؠ��EL����T����Dm\\�hK����3��G���JKc�AH�����f=��5%�l���pS�T�?e>�_O�9�lM;�?ҿ�v�`�ֽ������cOH&��S� ��mn�@�7ekr1��pe��L�� 7���M4	K^�Z��>��o~��Z�S�c?�x��®[0^>�����ՠ�9ݏ<Vq�)Zgff���������4����å����D@���i��>��%�l��a?;�Pm}=��+��wɎ�I�Ch쭋����1.[����{�D���Ԟ�>��/s���3K�������?��1=u��2�s�󻍕�.ݾ�>��]�������qq��|%����O���fp&R

�,��}˂q����{�5c<V�̛Ùfc֮��[W�v.�h�(N�����,,�$L�5������|���M�x]n�Xo?��I>J�5������-��҇�=���~��VX�H�O�lq�o�4,�?k���8@����l���(�cqt�g5�<X�pm�������g_�(V�hnbfe�:yL�������ir�̣���}����,��YLI��-��H0r���.���S.q����cY�� v�-= _]<p������B�z ���R@�ڸxl:F�!����醀�Z�R!���0���-���F(�U�rO8S%>X]�8��V� � mG`A�0հ��Y�'��/��������;շ������d�M���%{}u����a5�0������4��2F`.���N�[�JJux:�0�X�n@>�M�|��.hX�N=h�X��-�d"!�����6ud��3*��BS�v�sa�+'@U�P��5y�S�&�ZJI�������%�������n�����v܍j�eR��
	����ab``4�\�n����.[$��$	5���h_� ��t>[55����\HB��O��C�Y���$�b������b�6p!)Dk��ЍOs�����{߲#os�rڂ90^4.�T�^m�Ê$��R�J�7L�w�l�d�Lו��tY�n]�&�jqQ-+�~�ZG&����՚��Q�V^_J����!�pq�qH�{DF�j������I}*ҭz7��t₂P�����8��:�b�h�p�j��Hкޡ!���DF����,(}i[5�?�݆͑��E*�) ����vQ�Έy��hI]5k���/S�sJc��[�xJ�U�/�A~��,s��-L�i�;�F�ݩ������K6`��P�M�n6F�E<+���QC �A���Qi6�y���6 �����F~��I^���NI8 �K
**L�u��!^7�"�bu�I���	睋K���X���1�n-���j$kN����3ZV��_�n�V�y�����|�8Y#a�>~��@`��}�RS�b�?Z�(�����:Bo}��O�p&r~�Ohu���V��G�XZHj���immm[W6��ݽ<<<|����\ټ����'K���G���U��T����^ƞ(pg�L�L0ݫC6�B:(:H����K�j蔸a���у:z��$P�0C$�)�cra�c��"t�2����E`�Oٸp��ut�lq������V?��z��I晇�����Ò/_��x�g�ށ�s4�����$5H�Y�e�4mYZI�6szCDv+k�]�:��(��J�׍����ec���\���xK�nrխ����
]��tB���Zs@]-
(.`�7��� �J4ōZ��q����t�zhD���K@��3r��3��!���k>���I�th��w�T�[q
\p��|����N��f����(쭍MЈص�E���A4�M��d��Y��A��gs�-��߿}�FN��O.�,�0��$홌G�Qw���-h!'�|l.��)cʱ,�7�|����*�5�n�M�8@�⨅�UTTP�^;;siik#���zv�̔�m:� �i���lM��Ke�cI	쾥ȦÙ�8����c(l�+K>��5�9J:�����&��V8A��⭭�� =�4K��We ͘��e�~~
H��E��>~�hY��h�qy���Ш1�<9���oi�7������dWϧ��ݵ�^��t\�M��w��PN�5�{* h�����.�OfVkϟo�g%�F̮tE�l��s���^���$X���٧<8�=�D�s6�م�-��� 9��\_`�Ǵ ��1�w��M�F�� ��fәH�oǢ�إ�v�?�+to}Ƈ& G�U��4D�
2��;�������~���H+*Qoҹ�����̲N*HNU��� G�o��8��C+.$).�wu�:`���x�<��Kf1}�W���璒ps�;]7�3G�\i�����ce%��+�n�{{6V���@�`����x;ɚ('|~�J��j����@ )��Á�*(���؀�a�a��#v�sA Wg�����~\��7���r8�׷ұ��{&8�m���g�C�YF̌P�%E
Z��^,��!a����z�MO�$������͓Ό�.ƀ���U\쪰DoO��ǘ��o����[Z@Z���A�2}|����i��)�k�|{���������쑓V+g�-�(�T�K�4�u/��j��,�f�P�u��/Q�Ќ�=eM����������8�s��� ����lf2*E�ݎʫ|U��ٗĴ2���������c�Cr���J��������R�"�D��"������N9����67� R��r�%�-{Sg;8vFǫ1_o���dH@���ݩ������_����0i��69yy�#Yլŷ�$T�{5���D�z��	-F��>x�(.nԴ���v��h�ԕړc\��5�fLkO��~bK�����\�TIY��cH$�B��k�!qTV'�9,4/@�z@��������h�y�����˂�l�!�(B��}���BJN^��<Hς�/1rDa�Ҳ2��ˠ���Cf��.���v+����rf�cb�⏏���C����G�Χ�7!��,���`�7�AS��b���*�k8��ia��mw��(�FσR��ot�ѱ14��U#�_�����k"�5a�����!��X@DHX`UJO������il�M4�@m+�w�Ci|�`���>��������������Ņ���:~nd���H����F��<����!��ӗJ@��ht�CfQyo6|�<����� ��]��t�8I((<x��1�%|�Ͷ��|�l� K'��H�t��I(�-�	,�^uS68�n<��-����љŁ(����<�;A�����,���l���63[�FI��<� mE�Yp�����D�.u�[�uqz�1�	 �a �k��U��Q���;��]�^��rsy���;�����ㅑ di�M8iә�����:��DO���J���vMNM�1@nL��n�Y��@�i*煹s}����ڲ�C��o-�����-�1�_��b�~[��Bl�Ě�KG����aJ3l�������E��АH����5/.(���I�͑����>ќ!$\�f����-c[��3Nd����]�s�)��-Sv����Im嬆�"ܕ�;*}m��0���	(���zAAA�����M'}Z����=O�<["FVkc!)����O���۱{�3ј@P����������q�����v�zܙ�<��Ɂ >Z3
��0�q{S,{$����b��I	6�!��4H����s����C���o����fk��}�u^lE��!ہ���-RI�8�|rٱz����G>_[�u��	bO���u�(8�@\�%ft�^�00���:8���_��{�ü��cx~�%�|u����
N�	�9�&$"Zz	z�R��3�Gh��1e;fĘh(V�<����x�4�{�(�u��� �C0�ѥ%���6�G%������rr$1D=�_f��2�Pŀ��uzn�9����ȴ`��CI's:F���-��L��$r,�ET}D����xAT�s�4��]���ђh�k��y��GIt�K��L�{�E����㯧��&������-��gR�Խ:p8ꖝ�����寧��Ԝ�+�Z.!tH`JJ���5�⚩}w5!*���]]{v�.N��~_bիߛ�>$��2iY���~N��X)���Q�h�t��̽!������ӽ�C���[��q�ys�S�>�	Rg�=���Nl&:e�봫�2_�j�����P4j?U%%%^�����,��y&߱��@�H$�BƩ��@)�W�����?5�=�\��A�����[���SW�SiK��/4��P�;��Y;��c�o���� ���yP��wG޲wbd�,�K���JJ��lrJ�3G����B��2�ʋ��xz�$�<~���6��Z��vv����l:�����5c	9��+5�5�6C�YiKߑ�@���_��z��O=U��g.T[��F�g����#��7K��r2�(o=9N=JB��Eo��X��P9�m6����w�����S�����ë�]#�f2^/����|á�����1��j�_͖���k*/����,��B�?���V�y}�:��A��7ߍ�OFl:ա�^��O�{�c�V��w�+�������l��R�IW�HelW^���!���CP`�O��?�OGo���͗���Ѩ_ˈ�n����u������=�zL��8�8�7ͮ_�K
ec-S�t���[9K�TJȫ�={i����gf�I�k�z���6@�E�Bi�m>�8�C}}_�����D8�G̍�fJ�0����wvv�'��#M��X��Ie7����d��y+�F�hP��2K5��:�t�l-��AYKC�˳�@���k���p��4j;� �&}�U�H�'	h�h\IB�|�!U�kn�u��e�U���
�Qǝ*�k[XX�{��yQӂ�R��?��Q���~s��ќ���~��l�rή�8�P��%��l��.���o1����������ؼ�Z�4v��Q��� F�7���V$��8��Wk�p3����zp����߿�G��N3a\�)�|w���DF��i�����TW����P��;� 4�¨F����,��'�[�����G[���V�Uy�f\��`TQ^.f)����4�� ��?��݄E�~e)��:��'�HFh���`�nE��DD��l�Q�r-)�8�:Μ��y�f��[�6/}�SƢ��& H!��d�Pz֩X����_���@��)���'6��۳�N+��F�a�VZJ�������՗t�{�h�Z=c���Wcʗ*M0؛҂8s�S��ODt�̥�u�+�Р�<�S�4�q�O�������%�1�U������-��y�k~a����˞�ⵓ��DD��k����"����mWE�-������@=Y �����LE�3�Lү�� C6@��5�:^{�tw��n�*
͍��	3;\l�����&�Y$���D��Q̘�ؑ��󋧖�BF��g��<�6�����T�X�S�*ՙ�qe�<V�����" ��ip\r[q������I�;�7,��W<�l1�{���4�������T�%@���s@���r���{\�:Ć�y`�{�1�5�}���u$�k\�^W87���fL����!�8��٤���6t�9;u$m�<o��߭���)3s���Kh.K�Px�/8f���V�n��g�T���NLo����S� ��u�w���b�cu9������ͬ�����yy���E^O�zh!��*�#P�u����������Db�K�cӁ�%V�� `�5�	{K�����`-�>z�ش�2ϙaEn')�Wm�� ҈Y���=��e\�I�7C73DR�e?C�cx�!4�輺�����j����f���Ɵ�:aH�qbȯ���V�[JW�Q3��l����B��"�
a]T�^S`C�����V�z�G볋x�z�󴨨�Q���aB�p�n�=gv&��[�f��Ў���[kkk�� Ҏ	���׶}����fGe�x�&n�:xP�d�������ͬ�]0�lV�f��qM;�&�����F��?�<۝9��+����ē����c�LI��3v���2AƜP�RF'&�@x�f�U�==_�?���z�F��~�ZO���X���R�}(3	��]� >Hp�)�PL��o�g(}^�:}�I�$�C�A�>rrr�*��̷z�@��#�����@n�#�3T�Q��^7�;C]�u�{\���` ��!h_
 2�˥)ۍ�R�{j>���B���z��x�~����
���L�����TC[A��_����]&�|��ҊW����i���-}z`&[�S����e����r������5�6�p�s�c��V�A:8 ��åÂd��� lH�z¸.�8������p*�P��c|�������r�u�A��|'�J6C����� Z˂*�9�Ө������Ģ���^��B�͜m�k�&uh��Sw;I��*�$�3 l z���Jp�y�j���r�/~��,L-.�q�l����pTb-��ۇu��[�~�u�@�98.���,��	�|"�*�04�����+��� �%�XY��dv��5'������C�"�P�b'����,T�l��v��\���q��4`j_��%S��$:�$2V�6	�;	:�1_���l�'�x ��s�CM�u��7,�?���h���Fc�_�PZ�d>���sh��sls���11}*�9��ߟh#q��#�QqT���a�|`��Q�=�X�����F��N���E
H���)D��䔔z�+�� �������ʊ��ׇ2�������(�)���,�үa4��*ZX�玉S�mA�͟��.�M��]B%`}�k��B�,_�
�lE��_h�z.94T68Pק�?��}��-v;z�=A�Po?��\��ƅ C.����&C̨���I�8��U��Ȑ<.�:���vu����t�4H��x~xwp�M#�����ӧ��=!�����!ψvP'ƀ�(7hq�K�5Ru�ܚ!a����{�¨�t� ���a�0���S<Y�,�����P��;)I����8a>�4��m�cɏ]b�DM�h"..�ݰ�m�9�?t�~_m�m�}2^^^��F��?��x�n�&�]`��ȅe����?<��X4���>�L9�8q�8�y���%bS��Qlf��AN�>Kk� ��z������c���C��oo���;Jꉣ�Y�wO%''�c��Z�L 4N�a�z���z�k#������ps�(�b�QQP���D�A�[�{Z�z0Dz�%�h�iO�PN�D!�=�7�Ul!���Lt	�;G��$Y��Y_�� 2�7�^9�CjiբA؟���\GD/j1$~�q�:]`�3dccs�"|�gg��j4�xq��&��_���O�\_�}��B<+b�e��^� �H@��[)J	�!�P;`�Bn�#��<���n�2��[��hh8xuu��G6_QPRޛ�V��F[��J
C���,�|!�wu�K¤Z�l���%t��$�v ��]3p��;_+�+���p�^*�C}�{tc(�͸O�����G$I;`<\\n����Oq@Ș�%aoTT�����y���1i���B ���C?}O�{{�!1{�RjYY�8;+�)�����<������Ca�=Q�%�XT��OLA���
z "]�h�'�<j���:Q��u^2[`�o?.�����<Z���7�*H�S�E��1�x��d��e���w��j8YZcp�2y���C)�x��rAA�>yVs�w��VS�A�����"��y������AM�]�h�B���"EP� �"�H�����	%�J���"���Q���K�Dj%9�����?gμg�3�o!${��^�Z����PQ!���Xt诞7�
ԑ�WR��<W�������(~3��� X�m��� ��dtioR1��0��ˬ�Nb:z��Y�A�E�z>VȢ�BAn��4t'��VF S!�3�Rk=�_�& gIs����!u]>D�~~�/d�9&:�UNN�d��O���D���0�)�~AQ11�fG�m�>���}��wE]e�^X�7��/Sc�d
#n����=�AM�I&��T��̨C���Y�7�}�XI��݇���8�r�ox>Q�����a^��T���-���M\�ຒB��e�B#�ʆ��$=�&�v�2p��O����4���a��3a�S%\� ��������l=wirq�D7cF�~j�'����pZ��p
E �X<�S��9?����u��E"t>z���K��DM�=9����:LV�����~�� n���pӲK
�]�v9�ש��刢b4�i#\I����#쐻�?���#WG �>�꯽{��2h�Ү�/������'��ё*�	`ޗ3C9��v���
&�%�L�x,�k��tC�˗/�_+wsut���a��iR^�ɇo#Y*�7����k�&�z���.+-U��aH�zg-�F'������z��w�����)���S�(
��a�`������S�@V|�g*Ć|{��~I��e��-�xDC�> }%�-Jy`�A|e�������P/Yҽ-̌}��<$ґ(F�FK���OT?9K���l��ʅ�dw���TVV�H;�<�34LL�]:yU���8iюiV9�6�?y���@�N�;���[�&k�s��jIⷤ�hg��[��6fփ��nQ�lL{?+�sO���m�|`�`�>������WTlI-+)�\Y[�Q@�{�RZ|n~�H��&۫�{����Jw0-������	�1����7�����m���O�,�Y[� �'��:�/_i.KR�9�����՗w��&��7K@�:A�?�|�z��'nz[3:::`|�4Anp��i���W����ia��h�{
�c0n��~�`(���Nq�ij��Wl<�
̍'������?<l),�ko	�x�(�
�B� �c`:M�4ed'�������uq�Z��O;	��(@\����Ǫ�7�_��dR���{)a�թ�)�X E�qkk댼u�m@d��ō�՝�7Ww���M���b�J�g?�����6�$&�`ݍ����L�,�;M��ݼ�
:��ýLI�nkB�����9�5S�&&&\��JR]Tq~����}f)B}��H���H]W�8����F�P_�"�HYjj��߿o���qD)\�C�����g�d�x�x���BTDͥ-����.f_@���������"G�:~K��t�@,�Ib�`�A(�'�e}<��0�ddi�P�t�Qp��@���o��/���@o��MC���r���ia�c/��OӯF��}=�pÈ˞e1��]�̟v�1WCC����9�����|F����îx���e`��ѧn�
u�v�~������g�oIJ"̽��,���===�m�a�k�u�?��1t��G -�^ziH����w0��ggg���]��_zP5	���X� ���������w�|���U}�H�*�U�zX��gc��ڔ�]~jj�����FԈ������q��UK������h=ޘQP;�����7�Q<\�����K�U��7�>�2`SYe�,Y��|#��[v��V4qXOW����j���0�k�������Ґ�
ra��2����|L�0��|{���=*	~�r��v�$;y�|x7��KA�~9�W$�?"��?B��b>˿�����z���։�]�a�^�W��ž�Vgp��H_c��[A����?l�N��M"��d��ND:A�JS����z����"+F����hJ��{��+[��:HM�ĈS��p�C\*�r��,�ZԠF����cA�|y�Z�'�V~��&��l!PK�@���P33+R�Y#�8r�ӊQz��-]��� o��1��������Ld����^����,<�l mYv�-=ȥ��)~���Z����+$3485���x�Kk�_V���f��5O^J������A>����g`O�`��g�NT&�5�V���\�+&�z�#� �s�����١����w)�2�5Xi�����k=��O��?���AU�f���z��ޫ��L�N�'������b��]��q��ঃ[X���h�*��3-�f�QgE���|9�|��P[��R1í��v	(����Ȼ!U[�|HY�ô�dl#Ҙ�^��_��Io] ��t{�F��׎N,QG��d۬!9*fk�����n����1�ݦF{�;-��m�ւ ��M�"�(%�%-%�A�[n�L��-�w�%�5�L�dxr5+�˫��T�O�mQ�`�7�xb_�z���-�0��DL���Ъ�G��uE>$=����L��6��W�֌!J ��Q�ɥ�t/�Ù�t������Z6�)&Y+�E�z�.�l�&�qA����%�Д�# ^$�c@-��
�𵜗ZG�!YԴS_768��\,�.��u^@���Q����9������.w��&��։� K�)Se8O��[�`_Az�s�[5��y'�'s.�zSi_���S;>ǰ�>����^b��z#���፣�ה�V�" f�r��ڨ3 �|�9�5���ʫ�9�-�zqK|u7��'̤c��i���V�ϐ�����ü����n�P����<�-ߊA�,@�GX�BxQr�zg���vО�"�$�x�)��')�i��Og:����o��b����;�=��e����3�ɩ�.���gAd ��iJ�g�_��I\�d!�5`B�����}E"�#��
�K]v�(gc��u���@ډ]]�u�U^��}�u�b��/��f0b�ǣ�rA�Vn)nP3��eQL�G���?���ѧ}�G�9�r����	}��O�=V&��$�i�J�^r�Zφk�'�g��߫z��v_g�����${�b2p3Z���.��u��k��~Ӆ�OU2S����R��X��̵L�c�@}>5�6�����ģ�͚��e7?�
���\M�辰^��?��	�	6r��Z�RS�R��6��y�{�x6�E���*�8cYe9��%��8�U𤌥��x4s�+B)^�^2���,Vu���%����(-��BS�x*�Q��f,>H�&��<�����	N������(t&�iտ�O>�^1��M^N��WK��T+M��Q��~�:�#ِ��1,�³�J���Hy�Z�.��&�1���5��M]��h ������d�6LET,�Y���i�&DVr�}�K&�u�[�?��Y:���}��P�KR���D ��Et���)�5���k}�i�#(���Nt��-Gۡ�����f�D̍��Op�u�zL�"����p�&M�D�>��k|�/
��S�Π8�|�U�a�^|�Lj<1�Q����$�O]�	5Ѡ���[&,Q�1��jo^��`���|K�i&��z+��E�e$wa~���6-��!(j����vL��������*@� ����x�w]G.��G_���)L�(�.�P�U���D�����	K�%�x �m����ؚ�{���V�����dM�ʽ��d��o��v�R'���^+k�<搜������'S� %�V=g"�X����%{��2���Q0kK{5{��%R�Fc��oƦ�,ݬ������a��sUmU3�m��4^��x0��(���JQ
�3�-��B���Ѣ@'A��݉?ZKj��S8�$iu�
p�p�|	��R"��P�Ek(c(�)�������:�f�!�C��#85в����Zu�<2� &V� g���3@7F.JQ�*B�%�5e�+�~o{Y�_|�Z��[�,o���r�Ɯ�<�@�u.q�JotmT�_��$�Q�������&�p<�{�o�X�#������D�o ��,㳊o����Vʬ�Q(�(b���,�.�KIY���4<<�A�Xқg������d�M\ջ����<���=X��DY�����	�]���zO�}��N=�U��j����c�~�����e7�s��Z�ȼͥ����Se�p6q���\������*_o_x��wT�`7�0.�Mȃ"|�W��Y�#��/P�����y�Uỏ6\Rp�<�ro�Q*�,��5�%/���>2��>�EpPo�3����~*�1,���wK��b���S���=];��h^�<��]��������t�|�|�08q��hz/g����O�uV�aD�P����I�j$�������-#}#��8��q?<�l;]s�ynu����V�Y$�f��-N���Ꮔn���0��A�H�V�O��@�yw��:]*1����7��DP��
��6����<w�M���؅k�M������{��
�
3�7���i�D�ɫaYk#�Qq��R�ʨ���3�>}z}�ڎٓ¶y��(�|#>ĩ����S��6*-�D腖����M(��%�|���7g�=�Q�����Ǚ����>+�VVׁ���l>��}��ͅZ&頪-�,����V]e��pb'�M��͛g"�R�� ����.�lt~���Qw�2]��'��z��*�"��C{�:	����"(��bqح��������IY���g�Q���O��ɪn��>&��2"��	K�������n�,��4Y��drݶ�·i茊DW�ds��[ -�8VV˨�RK�w�!��S�M����m�2�v�nYbk��)�oD�����zm���z\���sp�F�~�)�Y�D���U�#O~��ȧ׮�3�N$�6;�2F횷�܌��ny����XQ���#V�84Y�S�Ǉ�Ĝ�S���m	�~�,,,._~��{��{>&.))��y26��=�Eb�e�����?�C�E1�#��ٳ>|�`E�+�����P�g�� `�����d��%���pFI��C���X�x�-mjjw�yP}�3���C+f�^w�V�c[c__�2������eͤ�}s2�p�ڪ41sfqޘk�ZL���]�u^�i�n�%��1��������q)��|�u��F��SB8���c5t�ʳ�%<2r������le�Ψ��jW�,'��Ix�Z�l�Mg��g?�y���ݩQ���u�a�%(�GF����G`R�E�};j����|��Y�!1�a�r��MF�Z�5I�� h0��Sl˞*f���������m�A�+e���T��n��t%��l.W���ׯŝ~��f:e�d���璤�����^���c-�:��|[�H����a9G�u]���t�
`&t(cU���`�H+^ ��@��l���n���nXu#�j�-�5MP��֫p�T�*���b��rCΌ[�d�ے&5-ms�Ϟ����X\6��Dk����˗mJ�&\�'\��~�|�&�+eV�,ɋ��:��g��|��g��k{Povk���}�2���.+�tٚ&�tQ��>r_5q!q}!�Q�A��ܳ�y8�9tu����i/짐�[��%��+�l�a(];-�J1�׺���D�h-w���ήO�����C<R68$d���z�y���/�̝��:��������x�l ����mjb�:;�o��ywo�`�a�ݛ2���⾻Nlw��:[0'bᑱp	�|\jj���F�Z�����#8�4GM��������28�35�(rx_�
g����bnS2��Q��/��U��%�<���Q�ZK�֘�8v�/�����w�|�k�~w�&"� �[�8���\� ��ML�_333wף�l����#��:Y���հ���Q����CE�.v5�!��9�'
***�ʞmb��Cf|��N+D�IXY�S9��O�KIn��]�8��Yr��k� U����i�F��wz��\�����O���@ږ8O�w_�>�B�F��VmlkS�;R���R�C>�\?��VY�s %�S�1�_�q��@:77gAh��@
�]G��t��F��FZ�����ugH���w��@*����ۇ}e�3Ma���fX�������6>t#���ٳZZZ�����"K5ٛ׮]�k_YYY&BQuSkVF3w�o��Gdđ��T^��- (P��AM��P9��/ ��ק	A(f�����%��-!��S�	y�*-�S"�,�<����,�W=%�M��s�����	2�G�i睕'��@�&K����&t	�38L��������Qw��Eo܀���/kW҃4��7��ث"l�*>�n҄!�� "������Mg[�ZJlM���^�O�M�ջ'��ӣx� �)���^;Q1�+W��ܦ�V� ���x���`���-�kf?�1��$Y�{lu��-�������a������kU��*|���:8zX��EZ-�)�\��+�l��Y(���3(Py�SU��~0���yVc`�D�w���#ώJ�=�k%�K�`�i�`��(�����ۛ�h2�r��O�������G���`:�I�b �WVVn�74�OAQ��Ύ�������[����.��ϟ_�����^&�(!�t �� 8�-YYN�w�-�t�47��������Z�q� �jj-��ROAw5v����YX\4��X��edd�.-�c!;00p���qe���S�'>Qc��#���@��/���X {M����B�]� O�W���Y'UŀПA�Xi���iC��߀t��G=V`�}�,�Y���|{��ļ�z�g����?{ju7H�3b!k}�O���;������׈*:�pv)��Z[	�߼k���%�̻x��sO�8���`j%�#yQ.l����	���ȸu�[������tmަ�����U����j�U)�|](2`�

�X�%���G�?8�4�B������S�P���zo��|xJ�%�` ��� �A�B__��wC�o�S���--��YBT�b<6%,@^)S�n����n���Pų�����h8���'����܄���A�ׯ_�����w������(d��z��>� �B��T�,����:Rb��Mry��e`��>	x��$���>�������\�ý�#̠���;-/���Z ��o@F@���ppqqi�W�[�ϧ:,#�3>>>.99BՏ�:�ֱ��2Vb�=q[Z��?H�*ɩ�$x����bC�f[>��������(�C8<$%2����g&t.,E������j�4_GOn�X���;c{>��9¡\�K�A�ҟ�i���X"��}D���� ӏRc:���M#����N�|�s,��1����ͻw��RRH=<`��c%q��o��
��f���e�{����l���%��}�!���|�;���pI���J�f��p�� �k A�y�N�������� �Y/��I �QGL��f3q�e�r
p�9k#�&`����k+�5�b��ٕ�m���c�^���m0ǇRR�6Rwy�&�t|u��ӏ+�>�3H��Sb�с�g��=j����������p�L��<4XB�oA���*��1��x�� P�[��,/_�\o�_��_o�1A��3b��̨ٔ��d�5�l��H>fO7@�ɩ��� k��f�.7\`�В�����1t��Q��5��Z��tݙ���¯_�.�4h���%$�x��1ϒ����ʲ�[���٨���߿C<��~F��m��rQev��R��I�Z�-~Q�2��X��ˀy>����o"�Tl?��^v��*��Z<�*"��kjz�v�IT�)(&����r's��z�.���B���K���%�c�z��.p�tJ��� t݀��Z>��h����'0���dN�kfh�Nn�m`����U�YYY�@���gL:�ip�+e�ˠ��x�����r�~`t9�����6�W��5�����,���*�x�.X�����]��sB��k)2��ǿ��eS���M+?��K�_�|���x�!��`�疻���\���Z>F�a>���:X�4t�IMy�ԋ!)��tu&��=.Z�MN�6�yƫ��g�	�	���Eؓvir�M�dC�ogK|j*���*-���=�N!S�q��_�}�be���k�J6��_|<�_�w}�n�˺o�ٵ��GEA���M�=���al�5�����1�~F��%�TRg���QN��F�3`j�IXJ��5�,��M)K�Vk��S���V�,�kų�B��]!�����\E��u-�����Vs�v���4�z�*�?L���T3:*�ZL���}������#��0h��Ѽ���u9]j0¡f|8B>�=>��llhʑ��R+H�^դ��n�*"�ɸ���m"���KCH�Z"tЈ鳆�!����R(��i#J�"*��z������)�Sn�?9 �Lz{=�4[��H�vx���t�;�/��4�^y�
v����ʢ�:�>$R�sI�����rE��ry|��kG��(�5Dv�VM'�<clЮ]�rk�U�J�W�)�����pҨ)���{��,��.�;,��hg0�Ց�Ю`0t�5���� �")�����%�dQx��)/Ϩaj��(0�@�a���hR7:	D�&f�R)#��<k��($�<� ����P��`='�����ރ����B���V?��P�.�Np�{^��K%�9ߢ�U���\��a:u@�v8�xP����1k_��-J���=C���t
����ѭ]����O��~������$��1��������
�Mo�����$N�V��Q�`���+��������.
.|��.m|m{t��d:_��}(�:+1��Bh��|@)�}��ϭj��+����G�8��F1� �$6�7�V|�~\�w�����;��l�'��+T�mOChMW�xe�}/�+$�+Xܒ���X���-����+�e���8!*5�s��OH�pA�O�צzoT���&WO��b��,M��^�YY�d^t��Mɖx1��s�-��R��O���%�|�z���?�Č�����x��N��Ô���k�
34��?u�cb���hG#ْw�J��q��l[YlE
@�_}��T��rjb��/��E�䊾��Jz��N�}N�u(M/7xo�%�D���Gkzy���Q����.��'�����O(���	<�I�_^�zYf0n��	^��a��5.�>�%G����u������{��/�+�%
=��tP#�ل�Q���FgZɀ�?i��)���p��1��_	�i���n�UOB��Gn3��"<��8{��?ޢ��0u܍+���&����:]7=ê�o��ײZ����'/i�*�&7�А|�ve��T��SR
1��f1�Y67X��� �gK�MbO J"N��Z��lFg��7�;̋��{��oZe�[��%�Z�W]w�ry-�E��Tt���|��g��(+%��mVF�r���V
`���F!���{��t���1�#f�:�}� �Mb��=	{�����ҏ�4�GZ(ٌ�c�]�S�v��a����2�o�Y0?j���[&3[(U?��ٝ��|֚��S,�Nވ*�)�w��k���ځ_��;�P��R�_�����ڥ��\=��۴�h���-��Y06����Jgx�eo���V��	>X=���1tЄ�ui��2H@h�O���{���\q����?~�osg��/?�MR"nm��#�wv��z��9>�Pb�ܻC�#���O�sl�V���;�N��=ZR��:��Б�5�5��%H#S���Y���ԈJ�*�[�5�S�;_<Y���Zz8c�Z�"d61:*�~H���.�����e���xD�2֌.p5L����0,Af��a��M����鉛�M��9'����t:T#�4�O�1�Τ��~Z*JE_�3�O��gK,3�E&Uw�!Mxf��<ig弝kd�pG<�o.�N/�f�rM�Yv�"���o�4�J�a҂b���Bin�_6���lNf��Y�@66�9[��}O�{��N�`�m��y��5x@�e�v�A���&c��b)OUq^v?9��^U�g�ev<z�)��Τl"���}����Q}g�c���<Kr���m�[R��_]�U6S|I��pI=�G+z�d���M���0���2��\���R#�~I�c��n�.���k��O��W
����l�	�x�H� [�|�d�-��G�)���|���XG�m�����`��xY-�ΩW>����|L��?ó��j��x��hwu�j��T|���k6�cwU����P������'$Z⋓D�GǸ�N=أ��w�]����/E��]�A�a,��b��Kzx�'n��I=A�K�����m���f*V��94��_Y�Yg� �	�0�5�}��x��٫T�ܹ_�ψ�s��#�:6�E8�ȡ.����uٔ��Qs%O�܉��Lj�un
���Ϛ�F�"���<k��#�$<�e�_�c;�Ϥ{S�]��B���*�G�7%�"�����
1Ѹh�74�����A�]�5�Fn����a���:W��ҭ���S`~�ǮX�Z��Q�:��?�X^L����츌T_�ܢk*�!
Uf�|1�c���K�2�ىy���gm��c�VO��AES�^tb���U��+zW�ve�r�FW��duOetL1�ǂR��	���q����P6g�oX䀱	�`�\�@�+s�Z|�l��Z��*_`	_���l*͎ S娺��v��L�e�'���27H񫜞�5�>m>t���8�bt�lAǁ��ӕGe��6�>�Td�U��v5�V&W���[��u���T�f�BS7�|�]����P!���i`+XzB���˭�˓d���*�6c����}]���?�[��,7�nN
X��o��j��hw��g�P�s���՚j~������iL��0�E��·�?Z�`��S�R����Y�G���yMg�w�v��v����QJ{��uﾛ3k�ڭ_m$|�E��f���>�K?>�ni�3���W#�ۏ���������#���Y9ϰ����)�������������mT%�ޤOm�Z��Ҧ�����1�$����e��������OD9�S������&a�5�|��~�+�16M+���4S��Q�Ta�P�Ż�5T�0Uf�"���Z�����^W\��&i���'���GHּ널ʁ��Zw������[u�߇���ۂ6m9�<|�5T��BaM�x��U����͝��LB��\��=�FN����	8�\�1v��)Oj���~&_�J/[ ���r.G�d�b�cb(��"�Z���ƗЊ�`�> ��{:�Q�: �p_޿����=�>�@�|n�A����_f����Q��7w�C]ڙ�{���l���I�=��>(ʪ���𲔿h�L2�tZ�/gޓH�M}�Srӿ�T|��{�,����SMށB�O#D
v���6��W�dal���}�-���.�27����������Z�S��!�|�,��u�5����lN��ᛶ���a�<7���<��s�f�h�8��P�9������IU�Ә�6YU�_����4Z��2Ѓ�!�t&��}�f��׼Hǽ��~��"�l�_c/�\w`���U���KA�ny�~W;�=�4b����{�A��mп�8'�Ge[�A�'����448p�9k����2i�%G��DV�ײJ@�Q$}�H��励�����U�Q7Ҕsy�Vp.���u�Q�ʫۧ����F�M\�7rО����Դk��>ω,�?��{&������<&��9:�l��P~z��z�#�V�'�E�}���O�v";h=7�r��҄��Vn����J훒��U^��w?�A	��	&1��o�v�	X.p�y�H"�����&�.��ɦ��}���˦~�TUF��g�U�i�-u ^�#o�N���\�V>
|��7s�bPσ�t|o�8�ԯ�&�ӷ�Q&mL����ԏJP�:�!�>�>��i���̋=�����2��k�l�I���	-O?�HX�����w���T^O1d�ר|������&h1��"��}����S
�=�?l�@�谵���d��Y�}va�����"�w�|�-�=x�gIY����/��N7���Z�xQ�v�?o���O��Ӹ�ygZr�̕Ũ�j��*�J��nX΍�nL��5��1O;�BH�A��{������xa��:e�92���ߐ�c�u�M��TA���4�/��^�S8.�4G���ӓ�7���;���~5Rd-!����݊�֭xjG&�W�'NB�(�"c�����k�6NX�c�F�[t�h1�{�oMT���(e��V�;�������*1u'���uȢ2�y�h��>�v�G�d����E��j��e�I"31=�b�f��;s&a�e!t���[Fnα_&G���8��"����K��v]��#U�Y�Nv@gqI����-��	׾$T(M��-�	&���G�rE�Kۚ�r �4�WD�|���]�,�ņ{�)�M�q�^6��G�w��E�6�(�C�'�\}������rIv��O�nXݯ�Y��\r�������}�*����&M��H3zŸ!�����y�);��v�3�.�"o,�K ���^;� ����� 7��Ss�
��#�L�n�X8i���&M��V �XV�+�$��=����r1b�ZNn�\���u=�X���z�����(r�;�[�>�ܗ'��̟�[o,�G�>���֑��mn��������+í?��<v�ny���g����ӡT���O��sk�ϛ.4����vN-PK��d�d�|l��Ԝ$4.�P�3�1!�^�s�U�����`����l8�h;uPD	�w��.Pz3���}r���Tu�͝l�mEUZ?�6��Z'�|ʛ�x<��g��T�����g/�e��RH��(vt�a����*�(�:�����J�Y��[��v��6'"u���a���?��Bqm0E��,i��v~DnA�
��
@�=��ޚp�H�S�0�(�����t	��t6(�4�~la��V���h�mﺶ��+���l �gk�jX�*Bu-\2�k�k�_(��T��{��T��\���ȣ��9���e	����ҹɃ6�L޷t<�%�^e�z���H���ll���@J��8�v~?{�H�p���~i�E�l\_϶lVfv����|�&�S$�����K��P�wq�X�O��@�<���D���	��񕵇�O�3��}��r��)��i�t��L��7m�g��#Ο^~��v��.y�3��	�k�W�jj�?����#�����P��O뮥���1*{�.y�#��C�Y���j����LU,�1(��o�$��-*fiX*�����R��Ь��IN6������Ѕ~az���o�<�̞7l�2�[�qg�H��N��X%"��~��-N2q�&��{��!Di���C݃>ц��~�w�V�%��?q�i��2č$_�Z� @
cl�M�O����-hN��|M� �f�\
[����T���H��n]<OFV��k:&dQ7�����d4�lyr�� gBrb[t!VV<�n��LU-�� F39��C��nG� *����;�{��Bʠ+�xk9H�pڨ&|�K�Â����0k�&-��K
>�Y=����#1Ix�$�/����W~J�T���?��#&
7%����guЉ��~�����;�-c�.m�W�W:,�S�"�O��heY�}��ѝ�{|Ӣ�~ �o׷6X����{
�#�CZܖ��QM��%Gf��~<�X�\}M�O�]HM�Hp��m'�1m�/Yj��%?�6���][/ �?֊Z�=��2us��ʹ���̽r>�»N�7�D�u-���\��a���i;�p%�d�������5�W���u���uU�i�7U���t㳉��L}\���;��D��ҧ
�Dw���`�=	y��%Uٌ��c��\:h�ˇ,w��]�K)��-�]7����J����������>!K3;��Hu���v�1ǊyF��#����۞��o�IF&&I��͉���`�}�R�[n�-��%��;4y����l���"�*�傶�i؈���ƝIuz�����?�V%�.Q!���	0��ǨtͰ��=�0��@�k]���X�շ�E��ynR�w=f%�U�H��OkY�WcePZ�]�WtKed�׾�U�ǽ���)Z�#�-�H#ˮ�w��^x�߽s�����h�_��m�I����jD�����=C��}0��͕�/�1uX/n�$���⌥0yӆ�{�f"%�[[�+wZ@en��L�m�­m��T�	~�K�ܢU�z�G��N{z�kA��J���ػ5:o#����|�y�6��K�EW %�BqǇ��{H�Ȃ�>;����ҕ�2W	f�/J�p7ܤ?4G��c�4�Fݠ~���$��!N��舘�6:;�3#��(x]�7.�՘W�5+d�����n�s�L�}�♽��}�n+L��q���OPG� Ǿ�U�N�Eźt�E��I�΁�*:sx)#q�$V�8�Ö�?����T�F2iA��]�aXҳ���O����#�'A�a9���1h:�$�L5�M����W��=�uY��$Ұe����Gb7Adp��C"#�ʤ�Qӯ��r��ߩ����}==o=�S���*����5�~�kJ��	2�j�N��^F����x���%*��ˁ�ѰN��n���"�b��@�������
���p����ܸļJ��q쀠�\�p&$pڌf�7�_)p���t?���]��xb���b�����X�>W=�ѭ��6���쵍²hs��>W�o�ԥgs-c+�������c\��\S�V/��q�/^�|5�"�7���~>ʦ�F���"n��l�I���C�e<��j\�݋ikk4tt�^^���4?�?6�ε~`aeͭ*X=׃��̽�������AI{���^�����E�2���%�t������o�9G*��g�bX���C��[۽�E����o<�X�~������ 7U�A���d)̕��Ъ�f�[iBMPSc }�x�?��wN�l��K�N�Ol��t�UN������Y������	Գ]��9�/�췔AA3�M�&I=6��\�����*-�><r�X��E�����.UwOϲg_�N�k^~�~����o)~��O�	�ݝ]41��
����Z=�SYV���2j����D�ԓ���,_L�Dq�s���kF;&ƹ���׳����Bq�?���l�K�&��LϞ,���zg��=G��������C�I��C4@~yF��Ӎ1p���ZCo3���I��.�1o���7�7�+w�Ztn$Q�ˍyo�mPI��?:��tE;�
eMz?Qџak�\�C�)*���kY+��:��©�/��؞��()���l�ڢ��3�nL>��vU�-�ݫ��
�c��������\��?Ѷ��#��Q�/�ǣ����3�3��Fgm���گ� z���������W�;�SV۱�/IA�K��"�>�*���f�n��ճ�V��/����SC �Ѷ�r��.�Zq������Է�Q"�c�o��l�ݯ#�Z��we��4�����M�~�~O��JJ�#~��=�Qj��層7?2�u�x�����h�s�72��\[  �ہ ���@���
����:-���Ǿ���1t����M"�L�_����ݷ�<H���������gB����[��ѩ���ݯI�U���L2����4l�A{u��f(Ĝ��0y������H�lU�0�k羜��������G8s���/�%��?=���( �DII9V�ZYY9GK�:��Y^�3-ˍe/N���w6��Rgpq"����Rf+d����͎���q�Iu[��h���1A6�U�w��t�m�mI_�K�V���܇�KSt���Y��y���mɑ���6�8�F!vj�;���&Y����^�9�~�ǖ[ò�ي��,w6�b��v��\/���!�nPQ�&rQ(KC��R"��K�IF��q���y.��b>`����i
�D<C��Qgi�v�\��̊���)�)����ƫY�&(߽�>!���UI�d?l��/��F��*!�
�[�yz��G
.��"��޻��K�8z
�t۫�2~d�;#���W��_*��i��x^.)�{Ol���k��j�����f���aEqG9�燍��bl�vm���5�����|�ut�P]�/H��#Qʪ{��;��}r��F�V��
ldc��?��:V���ԮY����ٗ�6�3��L���dq�Sc1Rl��\���.֬��г��9�1w�RѬh�zA�����f,��N,M|��Vr�~����[=����织�6C*E��(T��W���~���Y��n���p���ۦ4`��0���;6Ϩ������,��z*�9H2�9������#�������x-�s���G2?�FY%{�����z��rF&&aQ�ku��${��w�����R>|���ÿ��Y����`?��.�	M�6&b�&�$��m�g��a����餽�Ż�����w�?�fx�9xh�VT���w%����!��[9>ݞ�g��=֞Hx�.�5M|S$ϰ����\�����b|����{({8/m���ݕr�m���@*쬀!�Q��� 7>�9������OC�6o�K*:�%oɘ䀵@&}�5m��I�O���0i4]��be��GQ��b�Z��9������@q�.�0	UN����t9�-���ChJD��9�;��������G`�U�ׯcުuO;,<��w������1`�Z(r,[����0���L���T�h���|�����fǅ�Մ�����=����,�t��>�e���C8'{_���/~�&���V����X L�'�Ĝ���2Qn�9[�~k�$⾇|d0�_h�-�S��uq� (mc�a�_:4���ӡ,Zbw��q����|;�\�gE�	��W�刲5�Z)������w%*܌'D�uVi���l70лg�+~���D��U*�k�s#�D�m5n8��t����b����b*�DZZ�[�0k�' �4���V7Y6�����թ��|"
�{ɩJi���Q���ꫣ�j��		I���.i����;.�! �� �������ݼ}�k�뷖�׽��ٳ�'f�:h���gA
!�`���`��ŮRϋ�B���?g^��:}Lv
����?׌�3�ٙ���ֱџт�jڸ�����x_6�	]���V}]A���Uq�S����s]�P���K�2�BK��*_����2�oi��2�g?��$r����&gf>��|�0_i�!*��0Ǯ>��ֽ}�@���=�o�^1�f�w9�˄��O�fۋ�4[E��	ʹ�#�J@�0>��]�t���x��:VHφeO�7=q-q�'n$uArGՠ�;�7��~gM�e\����&��A�l��*�[j�q7�[�7������@������> �&&&?���\\8m���aS��Oh*���-�;�}���ګLW�2���P&�>�MW�h��:����QHJJ�o����E��������`�T����pu�rf�Vw�%��cν�z�-n5Լ�>RqݗwDkU+��Α�m�
���+zp����E���-W�v�`���6NW�;)�;�6����o��i�z;���2��~"Q��_�	f8����Fs⨕���%r Q�jJe�%��+\���,��)�ٸ\Xn��Q�s�8u���P��/Fk$D��4�9~Q�f�Ka}�5��՛��L��S,X:c��u�~x-��fC�p�ч]VЩ�W��C�3@J���-#���/$�wv��&��<��)���'����Y�>��:-݅�ϝ�hr\�O��kʘ]$���]����`�[�-�,]�׷(� :������Nr=
�Vf����Z��Wu��8�#�H�(N���@�n�b��t��{f����'}7h 6.�~~(�v�H����B\wcy�ߺ�z����w�[��X���+Ot�K�m� ,֡�sY}�ZY`P���9��ZT?-��Dn��A��/�{Nl��E�=Ꝗ/���D���ޯH �qd��-1a}9��, e��.[�Z4��\Bȭm�"Y,[��8p�̫M8��k��x~�ҥ����t7U?Rk�,�NS���("*��0����f4���M�j��;_�V�blVR��J3c�l^���r�Q6��'�+hʘ���:��~Tu((���kso��{S�;G���c���<�Y���o�?-U�%\���&bшy��`p�
|)����\6��	�]��=���U�>�6ŵ͗N�+�u�	�x.MS�j�Qw^&�������#�	�C�$#q;?��IT�]׆- �����_to�6��|ut1��@ ��S8�b}�t�����	�UZ��s���l�~`#�q�v�iT8��v�J]�/��w�S]�s���ZE��/�A-���[��Z]�?[��n'�J1�[��$�U{�u�t��<l>�r����)N�E�1�-�"��j�����8${��k�w�c��~@�û�����f
������0266\�
}��F��F
��z�\r�;�_6����%{"Hf*G�����B�P:嬭KÉy����\�W\���x:�����.5��l+�KsѨ����8���9�'�rYF�)�qH�G�bG�Ƀ��N�s ��8�\�q\Z��,*�H�y��}�38[4�ߖ0g�	��ꪰ�Q��Y#55�)�L߳U[4�xj,[4N&����<w>�	Vl���¤�Xͷ�a���>B�r��ې�{<ջ�
`��-E��j2�ѱ��V��Y�6�,�Ie����h+���N��4o�\��(��4]{0�*M#~�Ҫ�g0>Ѣk���I#y�����I�E-Å�|����5��&\�u|
^����Z���4)���)7dI:B��@nב��x�����v5�ԫ�w2YB�~k��'z`GB@'&O���dZ�l���A],б����=��m]�@�f3+�f(!�a��){oϔs���
jA�%零6Ie���4oqNAm?욖#Z����@=s󺍈r����2��8<���ƌ�PKg��3Q=�s�da�.Oч��G���-؋�˙���vb`��6nX3d�E��M�pB�/��{��v�_����Z�$:���z
�c�k���Fprig�,o�'F�y(�y���O��¿�99�l-��>����Ikk�{��� [��ʲ��De&��u����r�e� ��ן�^vHrK���b���6]���2�+��~�I伤��|�bra�Ȁ��aX���1�Ԙ_M�
7���+�6�1\l����E��˓�P����&N��eDs�[�}BW!�z�a����[�y#�ks�|Ec��Ы�~(�j5��3�{�χ�gwx82M��/�@����<`
ŝp];-�<-�dQ���7��5�������ܶЯ���Fa��_ �oG�U�m�!Ł��:'���M�~���f(��2!ޱ����q����b��tQ�^F���+��U1j'J���:���q)(��;�� u傄ל���q��~���Ј�S�9'�iOV:i���p�}�>̌�:Z���h8n`,M���j���/v{ЛP8�͎�woT��1�o�("�#�6�t��Sj����x�� Iu��R!kwö�T�eU�.ai�g�r*�sr{��">W���j-?�睔E��������qnG�fwe�D��c�'���쏐+$�jP'��}k5U'M��9���f^���S� qS��	3����;�j����+P:�D�^N�3:O3 �ٷ�zi�����3�˴�p����#���&�γ�-P��xwO�UY���Ee/�)H��������j����~YdR�@�@����,"�C�+\6õ@
�ǉ��iz�:������?�ޔ^�}������y����o�w�!g�;�J�p����
�=���r�5��0�ζ,n����^��v���x��J��=��ы!g���@��c�Ȳ*].�CG�`XcLn�@ɸw��]V�T�i��zV�/1�='1��������/�	=�Hjh���|�7��`�s�ɂ�����N[cd�nksŨ#������[��A]W`c{�b6���QLA�Κ�W ��Ư!����\_��~�Wr6�X4o�������V�^*��s1�k]������]�` �b���U�b\�R�lU!]r^#������ےOn��7�^G��)wN�.�-:��"�*n=���Ϊ�}�ҹ�Ds�����e��y��z��5��'PP:a/Ԝ�RDu�[?W�Ν�v[b^�ѥ'�C�w�ާYo��Ov�*���>.�J�M�.i;|��賁�)����i��D��b9.5�����AY���
��a|	rX�&���`�rd
�NY��aW��x&v��e�����ӯk����t����f����H�y<���N~(����J7«���V}�l(j��@`���j����]o�R��h���d�6��ڪ��\G�� (ZaEQ���>[�V*��1!_��1Q,��Ղ���4�!s��,�D���X�QQ�c�Ub�a���~��,י���\�9,8��n�/�mfnIƠ������7?�[έ�o�nl��B�R�@��v	=K�7��2�L6#X��t����]�sX/[�_�::k��\�L��gc�P:�X����qy{��"DǺ^���Si�yH�!��r~�PN�GyX�?Ʀy>������zq~���sm!�o"Sn�;Ѽ9��N?�T�Y�ug��^M?�u�I�C�?��Ȓ_�@S`���G��>� �j��x%'��L۟b's�S��񊭙7��ːg�B��h�@��[�Y�]�,�Ѻwwq�i��b�$R}/�f)��H���)&�4O��i�Q��z�`͟��!�O�2���g@9�nFS�E����r%M����rK�qz�Z�T�f�µ�Wi �8��U ���E*Y*I���gG�!g
��`�+ege�rZ�l+�����Ub,�HT�����-������}9r��1G�L��qE�G_�N�6Z���;+{���Ji}=���?Ϥ�%���o�b�B���T�#��#-�E�v��uu�u��spqH�	$��]��M�����q̦g��΂~]9�BH3`����Ux�%�5c�G�w:��=^Y5[���Z[���e��jrj*���e��yn�T<��x���P���R���˕�����kI_��:��&:�[]	j~!k����yk��4 H)qpW!wkyj����-��-�����&NO$����"@������){1M�,���R̘>���q�`�I`��:��.�Wx��c�q#�;�����{��LvS�Ԋ;'[�͢*��X5�[���3����tb4�h9�ˌ�`X���;w��$��"0��UU�2�ܸ**�1,\��dW��<������sj2�gLlx u^����՞�c5���<.��[h[q�4�ܻ ���	�²���Z�f7WS��-v'q�"���sX�|}�@�>�dn.��jO�t����?L�DmE��>$c[b��@u	����5�����	&�38X��)�� �|ӹ��>wZ3T���O�*,I��jߵ���U?�~?���6ku^��6���w\��6�#K���O��v�p5h~�!�]�>��-�P��*N\�����xa`IjC���{qq��!߿$)��=�p6ǜ�����4;[�/]y���-Nˡ�@����<5���I�>�wW���ę�]�
k����������؃�b�G������4�a�έ��᠛`�.+{�c��ȝ�Ool�Y�M"�#�9s�e~
��m��T'�Ѐ�j�WT��.��)+G�����_a��OMMuU���k��Z��~j.�#���ƌ|=����J.��pX1~7��n�Ѝ;���#u򐕓
{\f�F {#D��U���hH�a�*�./��c�+�@�W���G`sZ|������ܺZR@@���{��îu�-|�P����h&X!�z�-�p�������-�pj�uۙ���D��C�z5�&dt��o��� ���,b�nF�љ-="8�D;���5��l��K���Г�]�0>{lI]�����'�i)s��/Јgl��}Ϡ��!�U��V���~i�p����q</���F���+^Qk���!m�+׏��2�;�t�� �ۊh>���i)�u�2rǻ,�/�2��b�m��5��m����e0܌������*��}��W�"�3��%`H��T��Ԍc��*�H�d�=7@4&f�4ܵ�;?�2X�^�P�1$TҒ�l��8) ��*U���\Ξz+���7�(f���JCe�4�&1.n��><.WmM��[��C�P���R7�(#�.�<�H�jW�I���r����M�B;[ۭl�RO��_�����s�w�	��Otn e�'N�w2&�����b�5��t\�������k���&g�1Kn��n"߭�& ��+��	���鍄����8�O��8��*��Z9М3��C�j����D3sM�������;����r��4]�l�����V�:2�����CrO5����Ԗ�%'ۏ�Ѻb`�]+,��OR����p\�2a��p�gXgpѴ$�7�2q@>�M���q�)~ugu+��d��=�K<V���[�쌅�9L!�)o����ɗ6��0�6�B���B��U�O%	Je���i.ogq}K<��@4d��vJd�o����K�������lD9����t���fb�B�S�8��oS�90X.�;�n�%�҆�7�o~!���h��o�\�-��Dٟ���ɜ�� ����:|�-g�k(���V�,.YȖ'�-��E���mY'mE�N��`�����z;���Fd����O�Q�vtg��7��ٿ7&*��*�r+-~���-��E� ۜ{�4�K�MD��W�r���_���x��$������N艣�B	$vk6��Vv,���1��j����FQ�vśۜV��&�����}�J?B�����dI!a���+�x���Bf�p���;���o��ߏ��&�m��'�a--�BAw8�[��D�A��:7e�u���'=t���a��Y')0л����� rͧ�;W�q��L��٠���5�2���­�ŪϨwI���6��>Ұ
U�z�+�v������#8n�o�۹�&π���D��� �N��q荩�6�71H_�����u��Y�_(C(�����/��̠���ߵ��{ ^`�\OZș�|���*�{\�.��ذ�J���x�s��ې39�Z KS�8�q��el�l;"���_��؆��>�:�0�Q���w'�C�;*�r0��_cF��Ӷ��H�ݟ4��+þ��`�ۭи����3R��e���}60%�2=��-�U@��Bhf��RvXeN��[�h� S���?��������60��&�ч���(��4�M�A:r�ŷa��9
���������,(���c���3�����3�|�,��чno��ԣ"\�{��d�+�/C�������l����������RX�n<�a�&�����Wqw�d��]�RrHv7`0���ZV���MUT�E��� ������t]2�0|EY�[�r�@?�4�]���*��(,�')��h����ۣ����f?Q��[��E%N��W��K��^��fF 'c����%����z�c�ß�׼;�h�����*���r�.�Z�1B�֫�&�ޮ|7�E�!
�A��AE,�?��n�B��P����V�q8z1"�~��冶�.ɥ�_W"9�#C�Jo�[өܘy�,LF�jucs��K*��lp�u�d�6�n�t3��6��|�wc��$���Q�5T�4s��7@#��P̸�hr޹m�����$y�4$�r'���*;bVnT�#6�|�7Zx��l��\A3�/�灊7Hf|��������U�8o�����Op�,9.H��n).��{3f�ƫ:h�PV�M����q\��b�U�p�/�lo��P��8	+�^-WߣL�~��t�!z)&�^N��˭wԾ�[�)���X#��_�B�m�:�&X�o�r�I=��}2ǧމ��lor�����NB�s�{#݇u+��E��������;	�
�U�����2�dFVݸ�R<�x��=M��m�1�)�{ʏ
t�㆔��h8��D�NJ���1V�(�߹�����>;�����h_T9{L]��"���BR�����3�vBNQ����q��h0����d�\��W����G�I�� '�b�9q�yk��5�_��|��~�T]�~�x�Ҁ�gb�l=�k_���-@����"VX�3���z�����D�#&���h�jY*B�Ġ%�	?�E��j@O�h?ǚ��8���m�`6�l`@�͡B�+�}�����<���f�Ƿ�t��kv4��A�h�H�������v�?
���6i.��Z(�K��.^P�B�������qC����=p$��|*���6/��y^Dx�ݍ��/���<� �t�߻7�Tk~�l���F�b�����#:ZE�x\Z��<	!���p0Cᮉ?xG��&.�[k����#y�g��?�hv��.bt&��S��̱@ƣ��ׂ�,R�S\�|X�7��W�G8?�P��e�:�����ƹ�̪Q��2��O̻&����q�(�gR�x�~�O�A&/�#�����s�-?s�p�F`䒘�p������:��=�?�Bvw=q�[ȗ&8�LY��y��f������Og=5�U�6Uv�h��6�7>��*�
��
F�����I��v'�i��twxB�v�V,�+�7&K���t�*P�NQ���k �W�u�DW���C63�EVȄ.W|���DX���_��h��H�x�f@#o�|Z]=�u6��A��H�?��|������89�Y+X�B�X~���0��V+���ri �rI�3�Rc�u����������$��Ƽ�Ƶ�$�v	C-r�+~3!���@[.�.��a�%��4��/p��;T%�::��fO�	�\x^�� >�ccF����@D���s��d�,����d�V��$�(#vu}i�)�E)��}�*PdL��~*����{-���Ћ��s������������a7����,gT@���<a��i�R_�l���R{s��#sM���t�8\0���0��1n;s𘯂W�d~�Y*_y^�
�6�YB��vnk�R/2��"d�P��7��ė�Y�S!�b���M��=P��|[}t&`��L*�ꚭ���	q(&Q�����d��]{�PB�U7�*��,��0O�{%s6�c�$	)K����B��RfGĂ�>�JG)^�b�������g�V�w��yA�_��(�=���\�t��Yz ��g�	������t����������N�/jZ �	끏!�X`��e{&���v<J�"Ll'�R�����>����X�G^�}����/L�`��xV��D��}�iWہ����5�E�GJ.$����zݔipܥ���h5��D�ap[\c9M���ao;�X��8�f���M��O �f�=U�U޽~Vʑ�cO�</2���)��_�h�uH�8*�	�R����/ރnd�*+�O�-��uoe�{� D���(��f��E���q�;r�uFJnL1A��-\0K^Z����\�����ܲ]�fނ��6����/u��D�uʦ��&]�ı�W��1i|���2�e���!Ce�a<��r:����ѝW~�ں���b��.��3dk7�6Ey��p2��=��I*�p/ ���A�k��v����??�ϴ����;�F8R�2�hh�e�>��6�����GbCfG.�B��Q��d67�	˃�Q!)�,�
N�EV�������UxRDS/���x9I;~������-Lp��4x^b���ʾ� Z(4(���Q��!�d�Ӑ�č���gꃖ���/��9M�޳���uq@��G̉ c"���/R_�X� �q��B.�_�-��^�.��v�1��:�˃�T]X�qd��Z�z�����,�~�adpz��\6��Z��t?[�k���t�y�c7�Y[��)�}�1��w�;��7DKA݆�,f�Կ{"��p��:I����U�2��s0"�Ieg���7�#[���e��'��9-՛�ff;����Ž��D�����@HÚ�,��\�������MB��%�$��y��jah�� M�*�]�g#F��n��ם�RSfr!��x\�R�ֶS9���6J@�x�^�^=s��_Px���l���8�7X#����~m�E���}�cM���������]W���k��Qw�5">I�d����VQ���t2y�U����8foC��s��XV���%����	��a4-?0������a���R�F�֍���ϊ�O>,:.�Z7c�\%��oA�<\X	��Ko��F����9B�/�!���`�x놾|�R�/S(D5����m]�&辮3l��Ê,"A�pT��zOoqTs���� v�#�(�i\� ��q@=8
��+S��K{x����g��1�����ѫhN�2�$
��ݝF���D@�m+8���nZ��R�4��-����w��Z�ۯ�g`�y�:Js/w��rdlUW���L�C�t���z�=�w� �"�z@� C'��r��&"�'wd9�H�t���V��%�bK��D�d�$���%d�̄LqNE�����(�����8��l�Ƌ������;���n}��[Ԏ\�֟A�YϬ�>�#&v�:�K-�T7��5�#�<�7�Y������-Da>����xW�j����ռ54��3'~�3��nf�
���M�����?|��r5P���;Mس��k��ȿ����HD�?y��?����v���J�� �
F;�0�������=�u��k,6�^�c��" 
o�L�=~$�5��Cp�g�-0��M�ScW"<?�ǧl8�r��G��Jm䏵_ܶ�l�v<O�$��s�(�_Ĵ6��&�@Q"xB灈Q�^&Ic{"ފ쩻>�1[�c����]�x����y�x��앐�����'l�~��6 ���R���\wT,�>s��h�w��&������$�tG��� ��1g�]�����6�����t��� ?�ґZ�4�W��_�b��L�7x.�O��H� B\�AO�k'��e ��� ���h{��6�<��L�F��2�oA�l�/O����64��&,<;���<a���!IW��Jҧ)^��h���5~��{��4p`���VgV=�����N�dc�K�#huP֬�f�3v7�C�Ж�>�6�;�ZE���q��\��v����
�ۮ՜��[}��?�\� ����,_���٬'����O�5��ϭpd=Gu�t."ʌ�+i�|�o����g�`�O����%f�W���She9"�yn�����t������5|�M�����B4xY��)L�ؕ��ytA��������0��`��\��r@�Yq�Q��0�lg<�Wp?��Γ��pj2�E���G�x��'�܂��<�t�ur�=��i�Q!fd��xiF�/P��K<xV[��:<�j����Y�qס�r�D|�u�򌘝�g�
(-��w���#����[	���S�V�����|z(��~����O8��Ĝ�[��@���&��eґ���*��s�F^+�Ӆ���9,��� ��������v%��ddlŠ�V|�K��8���4�.�Y��&�E3켻�`��La�9pDtj*f��@����]��0i~�T�L��ޢ=Q����C����tq�誵�u��Ċf|���͊���&A��|b�哺�t��v�����MM��V�ha`!kղ���t��}~se|�o��>A�/���Ć�e^xX9���3Zi�z.�Bw��_W"���;f��3�w��s��'��~Y���j�ʎ�yw<�	{}0R0�Z���҄=����'f�����M��9�װ u�;�������?�5<�*���	�4�!�d��{�}j=�daQ�ڢ;�k�7��M�.]1�-O����?�H�@�����y�${�Ǭ�0q�4Yq/�6�,o�>!hE�Y7?MCt�h&'������hD��1_r���T���L�y@delI��*�9 �4�v�3��LU�@D�d��9T��p�/S�H��fn�.·\�M:�M�/�g����É�pY�]���S�s�l{�㢥��e3㇔�#q�[E�ޢ2w��U�	�c�x8R��X�6�~`Ϯ;F��������B��	�g~�)|�q����B�)<!G�zO�L&A5ے+E����@�9�	?��j|cr]'p�e���^�6����?�Q0��+4��-h%�O\�sn����0�=���	!b�"
|�$�'�noMD\�0��ZJ�mUW��Y��)N�a( �7��_�!o�]���N�>��J�����򜌂���W�d��$��d���Ό����P̘�AQܸSV?߿@-(��_"��=�yP�Ϊ�~�?�/[�H �Ԟ��~�E�'2��l���}[�[^p��`�q�w�ϕT�6�WG��ס�
�{���0Gx�]���s����n�5�X`xl�>T� W�S����7pl�!j�.�þ<,�7�G~������i���s���P��Z
��7hF�Q�ǝ����*f#݃��m�#5�k^��2��qӟ��7g��R�K��ϳ]�ݖ���ի���oF��:9h��v�~~��OZ8<�U��LJ�*A+&v�����Z5���?�yt�&	9H�[?[sX/�M�\�D�e����+�}��#�ε�v�a�w�"��%���$Wݮ>�������k�{�����+�P�ho��`1��s�Ցl�}E�?��X��5�i�Jn��;|`]����ޝ��Q����L�4[]}=���.G���aݭU���oI�I�N����{[�el����E=�MX��O���8���j?�[�乏`/�����X~��������^O�^�]w��s�?����ZY�e��>5
ɣ�r�$T@2&Kk)�����N\�O�a������pM�0�~%A��v��9VA�Ŧ�!�S�Uޏ#��O�0B�J�PPB�_T���"��I�����<��y$�oXʟ�<��  L���6N0���w�֟����Y�o�l���G����V���«��v`�Lxg�Z�&��`B
�-�nI�F����**6��g�VH:l���Hx�a&�E�|�nC'}&̼�|�&�וt@��7���"�"�)��#�y����Ñ;I`�4g����=�$�*�&�MP"����a�zř�h��}/�o�Z�H�̓���[m~�y:0�j�L^�>�˅�."s����+��������;��nA�`�|��c�]=���O�ozY�:w��It�R�ñF���eK�!i�*�4i5.�26y=�uJo���-Ԍ��΂���h�&g�`��	u���?��g��ld�,^_�zrOk����j�*&���
i���1\�mE����nd�*�;�:�d���-�$�a�.['ܲ��Qj�cX4�C�~3&���?�аdx�J<a�Z_�?����O�HCi�^~<��~~=�]*����?�Vҫxf ʑ�,�)�R��	$�b<:��:$��Q��ep"h�s��
��bo���ǛJN5]��{co�^�р��;!]:IO�ig�`d
`�#'R�/7&[@��#�N�J~�t���&�u@=}YV�#��0��s`Bu�?8(��ƅ�A5Q���q�|��C��|u T�kDx�٦��a+d�;7���H��fBxT�=�)c;�׺��'����S�>B��Tc��������+b{6�*|���:���")R���5�o�*ctӡ�����,X�WgXBVb=�5WX���j���#ï�rv���B�@���IW�w�9R��&%g�,3�K�Z�QL�=�>��Aw粚��Hi�\�����[�����7��q��)������Oo~=���m�hF��>�� ���;�p��0�$�a�K�?Ӈ�.��n��ot��_N���x||��	9�L��eU��;	�ۀo4a-oGAh�pĵ��_�	�}���zLYPPho��^c��"�NIP���1Q�y�t����F�n>~�V�^��4#���B���r����?AeWg^��[9�Ђ4?�'#p�zDx�D�9� �I���{Rl��dw��Ikn}JA�kRfܡ���#5�I�v�?z�z̫�x�;�?�%��*	D�]�^���� U2��RX{S;�m����G�gS㊄�����}������@:�nn@斫�c�/b�c�����t9�ޣ���>�I��f�6������21����'����L�Q,T��{�p��4�n�/�QWX_�ݱ;�
:�_�'B6��u��)Ph(:H��~᝽(�(�,z[���˲?���dt|P����й�0?��A!�HŖjHI��d��E������m�cl?]X<R�':�:A���1�f6Z[���29�|�*������P��ܩ>���#
�y��KŨ\�["��_�w����� i�fU����M���vj��$��^xԪ�obc��A("��$����E[)�9�4<cX�gs���C��!���_��	�����0vA�4����br����V��V6 B`�Lǁ���'�,�7f�4��S��x"D��"�W��m���Iʾ��]�u��#�![�_�~��gY�$���Xyǃ�YpP��������E"���6S�M����e�#��=���W�[J(�Sd�9��L��`L��<;��ʡm�\��`3�s�
�}q�*:�@YnU����QTY҂�Lγ�{܀ʅ�a���?�)߮x.݇н�K�N>	� �����T5y�O���ݛ�#���&_��*Ţ��4�ն�3;|���#�A���w�WQ�g��X�A2�����;�}�[�����ăV���7�܍t*�����6��+-��N(�=�)9
=Zcc%e^s�x��]� ��6��6>g�����f���4A�9&�b���K��L2��H0+Zª�,,�f��;�^�k��*oM����p��T�9&|;z��2�Y�Z�H��z�ƞ��A|��s�&+Wh]Gk�Ll'E.5��]�-��yYn���30FV�̶�
2���C�F�]"zk����<������s����غu����~It�C�'@2AMU>xO��1_|�:-P�i�f����mp�1�ɂ$zr/���P��C
�jK�s�lvOk��y+�ۛÅ��ov�RROo�O?��p?.�֯����]��ȯ\����'��5y���G���Yuyͮ�.?U+~8�&��+��1�V�>�㜟j%�d�I�G�Ǽ��c��Z�rXN���R�K�aN���5⿫20Q���*��P �	��|�ł��������R�ό���W����|j2<�I� !-�f�ܧ��B�g5��^guz U�N3ڈ�	�f@�U�@pz��<w%������~p�@4�(�GW9���8G6�_�A�p!�w�)Oi.���u����������jn*�(��= ��n�٪��N��f�Ґ�Zq&'�����!�vez�4��|�}��"�شݱa�R�I�����t�d����a�ΣR�Ƥ�����-G�������m�^|�C�i�G蓲���o'U0�y�>��}}����.~ُ`�8� %<ᝃ���ҏ���HR<.�/v�G{t��h#�b5P
Q��2�"�7_�! !�IG�
���+�w�<�V������}P��yr;r��3^o���Y
ْ4�Jj�x�t�i��؍���e7��X��?o���F�Oc,�v�I^qG1QY���f�m����V
�x�:X����5y�_��P>5^<��7u�|�4�CK�ɍ�}�Ȝ踉�<P)>�̘i�Sã���y��o��.���S��e��<֍�j�խ�-�eQUb�p=��&MҔ�^��⥽r��m�
:P!Z��8Q��>j���I9dX$��HY�A戕(>��_D��sAt5:bۆZ=)�1$���
T0Z����l��>?�I17�itE� ���sE�RZ.G�Vy�j<��`c6���f���XX��֫��4���e����ӵ����\�U\����[���1�����n����n�X���G6�l��]2o?�d)�doUǔ_ ���Jc���.��I+HLG'���:Pά;с�)OVGwm�!�۝�N���!�v��d�	}�Ӽ���+�)���`�<Rn�h��}�Z��{��0�/k�b���2�\��5�xk�.�ϵ�B�c�U'��tyaά������g�@���z��C��5�ڱ��16��C�2�G@����ߙ�E?0��������$�U
����I�fR�����<;)x�iEV�@Z��kZ��@=M;�Bw(�A!Q�AQp�N�sz2ɇۉ�'���|����nB�[�Ah�#J��L�����
�7R	����L�ȅ�D��ޛ^s&�5���J������`�M�������M��i�g�x�=��<�ț��t�|uW/��w�K4D�F�D�־���̐�W_��;��M���s���-�!�F�[?#��]���9���g�d���ȿr��m{i�Y.��T�����|�Z����t-N���מ�k����MD��{�]	��F�<�W���d�r9�{>�fjr&~���R��OC�Lr�[t-Oi���/0G������0 ��P��{�h,x�D�{� ����Q�����p3S�/"3�r k��L��z�B��.�Uu��;����8�G�:��y�-ȍY;��:���{N���� s�ݯ�=$�;쳄aGĄA�K$�&��M��Cv�B�-?jJ���I#�׏�<j�����n�<T���mq��2XL��.���e�-H�CږQ�ZֶV��庀�������AS�ˋ���2ôrW=>@��π%<��a7׿�}�X�T��t�	�<7m@}�t],�so�,�z��Z��=s�~Ė%�yFwU��i�~~KK᫿�F��pq''m�M'���aF�y �>����xla8����a�ՇNtݬ�?�y�)l��9U��q8�4M�n(���Oj�����2{��Y|��ޤs$Nᛒ�M�bd�]TW:b;	�Hm-��"�F���TCЮ(�}Zh�w��Ҧ�� \����}�i`g2�����{���c.l�Շ,V���*6r�����:��x=��������K�R|������\ˏ��t�:ĩ���݇T�m�;���2�3h'഍Ml_
���{���(ˆN�k�+�R�[��k��g+ Z��{���v4��w=�_v5�mۅ�lNp�GG�)��t��vwo�Ą�V9���R�.�؎�������^�#fe�^���"�m���ɪ�Ƕ����Y.��0"�7�k�67��v���a҈�`�Ϲ)uiD	(�2)T��m[��V��?	a�T���� a/��c1���ރl���!���-�14�Op����%�4r1�b2$" ��#Ð�=틝�N������8P�̋���!�I��:Z�S������kU���D�Zz���� ������58��J����'N둫IYʟR���uG�>4�ͦ k��@��{pe��:"\?���J�3`�cG
p|�Kc�s�6�ъv��P�Q����)�h�����l�o?c|Y�jv�l��;LC�ir��Q��8��'�L0	?
H�����0SW���2��%�E��6Y���šd�W+7M�r9b��_�����H:}GOf��NI?B�ٯ��G^���Y�O�Ҷo���X��:4�UF�������}uP\��� �@��,���\�!h�����Hp� �]w�g� ���m���}���������UM��{�O�>�9�ӷk���,�����M�b��Ӹ������d�S��6ki�k��lVh[���D�t���Nbp����2o���| q+��=���_�~�̌��Z�=�����e}�iY�E"�kh!q`tS����0��h�*:t&"a{޲pb:>�|�~˃�pM�0!%�y��5$�5V/����i�4r�^��3d���엡���̘���Svo���n��$�ѓ���l;���um��&��q`�|.b��lo��s�(� ���۸�*IF��2=�.�<w�㟃�Ҽeuop�i+��{5����>��PO}>Zp�.]�{����rhKYn��H~��_�l��yt�	(��'f��`Gr��2GԆ\@�}	�~�{ο�U��@ ��Fw����)�~�/�p���_ "�+w7�ћZn�:�E�iA��^F�5q3 �����B�ګ�E˨��Z���
^JL����|Q�n�3��0�-��I����h2n��*�#z��/�L�0&!9��u5��|��x��S����E�`jY��$s�%���L����j�=���G��9;?c��ײ��#����Q���1c�F7�;bHF�����b��	o9��T"/��!���q��P�������g�Z,Cͺ�f�°���b�Yp\a{��/Y��CW-���Z�]=��#`2�rA��/���it�@�Cn},��)��b���ݳYϵ��K�/��V�Q�*�E7�����w"��bx!U���Y�k���|���W�]"�u�T+n���d�'3�`#��#��<Y5&���@�a�V������(�u���9ϾI}@�0V��{v�r!�<u��
�X�	�����tB�jf�@sFqsg�rm�\�6��3Hq6��0��zs�}s=�6��v��%������z|w�4O�a��#�%u����tP�������ї(1�w�޲�i<UWW�t�"}��5��`2����}�T���|M�yH�_B^�/��G�"L�\��钂��E��@U�8�6�쬝1�������2��1��R�d��=;C�fn�FEo�0žMf>��>�0�����ȶ�]��'[���?�ݏ��=to�� y�����Ǆ�݋��$����+��\��@.�Q}b��Sq.�t����  �	,��� R=��!���1W	8��B=(ȗ����Cw�MSz��TW-r�B̰������F�Q�mV���{�c/���b�.ǹ�7?�A�
�w_�<6k-�m��,��:CdF%XߎN���t���qzɒ�4x�q�~�]s�"\>�QH |"�<ڐ-j�y�f �����"Tט��d�%�\��m�j�ؿ�� ��ku�f:�i��>�!۱�rQ��|#��z�����(���3I�<�[�,h�*#��F!�<c>����
㥒��xw.Y=�zFҝ���]� ��;���� �`����&Q����ql�v;B/�H	}�]�}�ؽ�! ��S++C��[y��H����D�����R��k��M#���)�,K���7p��F}Su����}ڭ����K�CPF)o��e��'��B>:�Vs��umXg̍�{֐(�<QW��L�^Q:����o�AD1��L~�.���FF=���yYc����W¡�����~��Q�}��b?��gR`/�H{@�1�K����O/zh���������8�Q�5,��$w��B\�и����M�+dG�7�ӯ���f\	x[�mc�$F����2^���T����q��0|m���I�^�l{��C��r�ƅ<vcᅂ��R����گ������]K�kd�}�kX�U5�tq� _����w��@c<]���+|�
��;zF���e�[���d$\!H<���)���a�W�q&!G5����G�n�0P�c}����_
	��z���4xЮm�ȜZϔ �u���4��z�"���(���H�o����,뷯3>�1"v�}��An	�O�??�l@%���-�^̬Q&5}��֏JF�<��,���ݍ�>�ag��ݩ�hi���
�=۵ȗ)�3�L9�l��9��g3�JfS-hS���i"��D��w_���F+���|���5*����F��/����m��Lu����9��#�Z;_!���I��W@��;���ɇ�.�ծ�\n	ڿ�:^Q�u$�H�lxLr�u(�����e���ϼk[�$���s	�M�'��TtOh�u���]�k*����#'���]�P��0e�1
�l��ǹ-�t͎���h�����ϓ�ׂ����"��<���@�����6&%a_[+�8V�ݸ;��yr�����϶|a��k�m$��F%#8�6II釓X���S�=e��7�L���O�'O:x�
Z�s��o"�<x���Pd�0�������67&�m����a.J���%Yc����XH�k�.[*�H�y�P��[ِ9��!�n�	�3�Q��^��G\�� ���!?D���"��1FQ��5�>��,���E'U�oױ�	G�HjJ�צ�d�(�"I�K�|�L#� &�4�#�F!� ��S��1�~4��h�P�Y�o����ŋ��T]E<�j���� !��������{�9�гLK"�:II!RW�iڌ�ց���)���}����Y(5Jܮ��;)E��؛�7j��ɻcAV�qH���Q<;���ݲ0�T���܊tI�s:�5��c
R���֋[;����4Oa�ň��43� ����ත�ӏ��ۼ�����,OXD� _�Z>�f��$�T�SX�h�|�;#sn��#�]Ё�ΏB��9��$�9��^�H���'��Jί�\_q�� ��h����\|Dy�F8|�@��n�3:�Z�A֋q�N�G�!�|�����PSt��5c�XYʐ�c\r�6�����7T�Ok�,��R^�'2x�O0U���v�1�Oy5�o��P���tLb2T����\L��6Az�����"��?X.�!���E�2^[DL�K���§A|�'k�f�:���\/�
�m�P����ڽ_$<�*��}�&]y��td��A�h�f�c�˚-��z�D-:5D�u-s�pa��߳��HO:9'��j��~\Z\1����M`f"������ZD�اT� �6#~���I��9� �s�+E���ƽ����N/�s�d��y!��,�R��8�$��-I���h�埿Ĝv�%��s|G"۬ �nt�c�ap�)��-���O�A��è��Ǹ�'����lR.cFو#����]�#��l������*G��������bO|�9����鱲ӿΜ��[�pb�=�l0+�q�R��MyU̵��A�,a�og��,����Ј8j����j
�^R�o��uq%���\��tWLM!M��sV�ar!0S�\�������HH>�Zl��e����=���Y�ǘjB��I�c�螣�l������>3�C��a~��tP&����|�U�ĸ�"����j�6$�x���~��7b_v����C;ơl9vC+��Ga|�����a�����n�0����ކ�X��yD���h�����g�Z�b�Oq0k�F�z�U	�n�U�k� "
�!]��v������ټp{�ď���"l���rr��L�� \\[#����;x�� �%k�1 ;"�>�O�|�'h��|�刻�5���o�}v"�,�RB��j��� )_;3��ʆ�eC��6eN�|�I�^�m�~� @�>����Z0���L	)b�}��=�×���TR^��7 )�d�ѼP=�l>,dˏ<�?��W?�$�>�7���?����Bn� ����,�z���Z���u�H\=U<�߇���c?��uܸ�?&k.m>�����_�$��@���R��O��� �eT6e bTU����2Q[1�M��y��ӷK>�� �Ԍ�i��I|R��c.TC���__�*��X�yX��9�&9��!6���-��l��s����rd��7�Wc玠�qe)#��7k���t���o\��l�Е�3�&xV�_s��u�%;&GI�.�@���c��}���EZ.���.����
�<�ā��5���!�ySн�peI� ���D�Y�:ą��� |*$�3�e8s�4���l�ț�K�Y6�@�7$�^6�I�$s(�	>@��}��0�4Vٺ�|�o���� �{����$�l.sj|*FbN�a�HaPm���Џ(��3t|t�"���,1�ow�MRN�*�0Q�Iu)�;dl[�J'�'�k�k607sw��<`�t�K/%���+�E}�������[J��� �B�ͫ��ӿ��߂Y�O������3���prLXs4�X��Q�����5VB #�䤖@x�{r���)�r(����am��W��F�\&�$�����]W��ݿ����D�$z+��������uƯF�ۮ�K�(����^�{s�l��Ǩ��u,;�ˉ�j���]�@-|�^����=l�9���v"�,Sl��C�����D����� ����Qkҳ�`�ʏ�,F�~�����FA\�VK'�3�ԼK���%P��A�A�l¦=�jf�g)*v�{�#������QU�
8�w��c��a���{V�%P��(�Qe��$uU��d���R�����|�����. ��x�X�' y���k�Hցtp��ˌ�'����p�|̵��#����<Z������˰d����}䠌�8V3n�!H���hGM�2���27�#h��#V���on�a,h��jx�>�\\��9G���3�r�԰z�� ��=�_�����K�ӹ�t�N�=Q#���;�?ta��_s�����T�+L�8~?U�4N�1�f�H-x3��H�����G��B���i��b�/��P�r�"O�IOUI�`�-�S�Dv:	O�^=~4���?mp5�������G��BA]D��3������4FY���$"W<�l֖�TQڬ���~�m��<�W�uԫܵ�9ֲ.����\�$ys�a.&�d�h}{v�w?Z�s���:ь���7��)t�wٌOɱ�myɢ v?x�t���O0��*��_���cި�l��x!ٛE�%�4d{�y«����u�(ZT!�W	A�^Ѫ�[��;�?Y��kj"�#��7Ğ�އ�:���1��o�j���������%V��}��Ml
���<�㌕���2.�J�M1?Vo9'�a����C�j����)^5��5�D?�F"G�c	Se�F��t��*6�[�Y�7�>�/锨GzN��%�!�Q�lB,��VYz��Z�V\�ŭ��O=F�>%ƣN��o0n|^������u��s����G]�����2u_2��Ͻ��J��A�\3slydX[�Z�B��<<�5�~v%VQ]��%�:�+�e��|�T�:<GLC<AT$�'rzП�h�M�̧[f�e3����DO������
(8��v��TWy��k7̓JҲB�ݡ�D@�C�V�]��X�p����|�M��$�/�u7���9��J��M�~KWm���H*�z��e��2���2Y� ����� �~�Y��vj�R	$�ur�3��_�J��~���<:� �G��c�40�j����4X�c��y����z^�!�Y�1I����ɱ�HQO_��j�����bm��i��$�Qܘ,h��l�c�ss�s�d7n\}�)$�z�!���k_4YL�f�����h�g�
~[�F}���H��� %�<��§ˇ9�	����e��͞[��t��3�'���J��N�'�\!�l�����J��1�{.{�Ѕ�tbL�;��b��?$V>a����=�<a+�:�|p#���(s���X,�e#��x��LIs�ni�b�����F�'�����G,<��1�R�'cZɕH�u祪����q|�h���c8=������`Uc#qt�v,R@t�dj̾�ygb�Bp��:�N4�kjCW&k�b�l且����,.E��o�{,\]J ���})OZ���j�`ZS]
;�����˘ve�l����8�#���
Mnd]WUGbm�qe9�4s�]�H~�>:�:Xs���|,)l#;m'���p�g�����V9Ä6;I�d*�r�}�CL��No����_ʵ�bt�@g�b=b��lNn�!�S>r���]�C�5|�-� ��6���e>R6�m���t����І�S*��lG�J������9���w+�h���-4�jYQ��r6��Ao�������81|z9v���[U����f��yW-[W�uu�'��=��������6�� m��-ɀ T����J/V�W8��P^-��H*Ӄv��=�Pwf�{Q���F��X#�S��Xs�����F�U>��Q���|�Y��g�H�#R+�^��+Ħv�H|�]���+D��.��4mY�t� i7�(m��_}�jia
v>#]`��EJ\h���c&�կ���Ӌ��ST��Q緟����޻1�Q�C�er��-�io�@�����^�k�Rʧ�	�:t]�'pz �t\��Ќ�X��Am�P@��4v-{��:J���r��1%/J�UF�薌�U�T�0>�����8����GLu�h˨��k8��q{	^�͓6djr�I���_�=�Lx�p���i�7��F�Iv��b,ݾ�����H��ԕr�4s��X��V�����6/1)X���5a�ALӚ��n�HX��D�9v�b����}`�hf|���6�Pb��Sί��#�IR����7���^T�Za-d'�7ޔ�D�Pr1c��5�>Z��4h�HciҊ���:!NV7�n���bT)�0����.���	���P�pٗ�^
!ڃ��}�_oȝ_��j��qmӗ��� �J�:S\6e���n���j.d-~�'8�D�{�כ�IϪ2J��h�M!�C�.��t�;a�,������R�aHY�����	:��5�y���;��))�D7�\�8��/n��c�)L��z'����©(�W����c�g(gn"�J�&ڶ]ZFO����${�_E���\	cz}��v�p����u^�7 ҺA�"�_�B���*΍�t=��؈��H��U�%^��������a؍�kT�a#F�e5�-�U��Ϝ�� �����pz���6]T}�;�M3&�R��8�r��ю^�",� ����J+�1���4,��ňȝ���}�g�(%C�-N��^����Qҧ��Z�X=��Q���2|M�.�'�d��Ӻ�6��T��И��3kJqqh�J9�� B9�ƛ�]�F� x0k�)����z�5ZG��@��������%�F(ӟ���괊b�#ڬ6�"d.e��w_�Ҡ�-��_�d��}��� ��>i&�Q����8�V�F���d��_3	����vA���&���ۆ�wD�&��_�˸l˽�px�$��U� �d��d�"��3��u���D��j�"���[��˟�y�rE���(�6�	J��{&=��1F��q�V��c�DůT۫��st���4I��Ih�ؘ���LT����C4e1�gN l����,� J|������� �&_�Do=�,�0B�j}�VƝ,�`y�����X��[�ݩ��Q4�$��=�9�S��%����;`��6��y���4��܎k㥛q�+���D���������wH/�����FZ2u�\�8�(��+�<a���>��wkz�]�|�24�P2��ɴS~�n��{{
��J!,�|��-��"}���>���pA�nS�q���?�B.���;����?�Ѱpr$��L����*Fi���ѵ&51$�	pY�ܵ԰�I1��e�5�5�meƖE�	��U��̯j�`��v\>��ʡ��%-�y�����ohl*I��~���񮙴>�Iw�z�@�jO���y��6Ќ����h��L^���un�YkO�;�u\�z���/)�.����v��	��&�v >�^2��ܫ��
�ۚ��y`z��3��ZJ��`ع�p�lC��7[���4OY�lC���|Z�Y���̴��n��?Rvm<|�M��:�x3n��V�E�|C�g�zK;��r�<��wB����y����LԒ楱�D�˿�T)]K|ܶpma��}�U�Wf��350�0��~.Fu����^�Zg��[z�R���T|���l�~�P��%k��:֟�`$:<��JU_5��qP���!g^^�d]�^ټ7PH�6u�E�=�"��{=�	�9�<�+���:��u\�pr�Yw\
s��*+}�8zd�Au8���w�圳V��Qr�}���	�裣�@����vt���jۜM�����j���i��~�2�<��S�^6����;�m�1�X��|��L� my�a�2>n٫` �~����Ί�-*������
�l�a (S}�Bo�R��k�xN�k�h�m���-.��LK���S4�-��Ĉ�'����>q_WY�~�ǑC�c��3O�����u:N�� ��,�B�'��G�ۄY��fޕ�b��I����M�p�����N�����F7�����n9�mY���
�g4%59��T�# ���¨/_l�[f)/�?rEm#+�Ve]G����we��IFyP�Q$� ����p>���ŸP��X�F�����h[��ca�M�
�tٚ���J���D�? /θ�+� XW�2�l�o�:�A���*��m/㗦:[����HEEE}�����I]@��򍍩eZ��L��݌]VD���>0���!�������d�SA���3?V ���f�к8k�(�z� 4�� ��Mc؛��!f^i��큓�d�tn}T��Ҍc�<\����:�0-�D��H:�\�%柹=P%%�9�n�F�YZ�(�F��Z�ݷ^d﵄5x(ʂ����G[�9�ֿ�,���{����n�m��,�j!Ro��W �������X��3cKxy��(���=����L��Mɤ�w�x�?�!�@�Ρ(��m�T�^eL"�]d�G��6�xI!���8Ջ���>�����{��r�, <��@myi�Y:@	
����y"�ܯ�~���E��=�����y�غ+le���|��1�?VZj=N�lڕ�J�v�T��9�_6}_č����e�9��HlۯS����g��{���Fa;At��;�r�+�{K�QtG��H��v,��D�P��{�O{�Z��%�ޔ�9-��"o!3������\���	󖥽i���Ӌ��xN"u��}x/�$�2�<�2�D3�u�''����!�k�V�X�V�WB �*nup�\W�����89-�N�"ô����nZRE�I����}4e�*���;R�"��-x�[��Alm@l���OGL/v�5}�H��K��XY��Q��s[W�¼�����ڒ���ӳx��Ṥ�M0�(y��j���}�´G ��W��k�J1{�)���{�`]��E�ā�_I�m�ź4�@��p<��ɓZ���ɕ������`,�<�d �"Z�)����E6v%�rޜ�L�\�} Q���]!0ͱ�B+��2-��X��1���u���"��6Z�($�T�;����t�߭|_�N����i$�3��O�zRƙ�@"J�ħ~�h=�g3h��0�Q%NZ�Y~���<����E���WEo���a��`����IZ�>��m��dQa��EF_�[ L\�{���5���X��-Z剁cf��L�B2�y��S����we*��޺��9\\�A3�z���P�Q��6=�͗�ע99a6�2�K�<�̿��4Íci]��x?4;{$'�g�2���������4r�en�m�]3��8����Ȱ�j�x:.�L:y��	\�4���)@��±��p���v>�ϙm�Y�%5� S�i��]=e��-�*V@����!�{Q=*�_��5�mґ����P9:.Ňپl�q�>�Rp�8�t<�y�	M6vNh�G�~4�4Q+J����a���;�6w�_+�W������;2uM�\(�q���D�w���p,_ķ��f�ג��Q(֔uϚ���3�>��x��	�R@�����.�i��զ����W(ߧ�E�\V)0A�׳�r%yP�1 W�D֘�Tg.�L_O3i��R�~%����æ��mڤ���T�˚�}� ��ѠOPv���Oo-�0�"��g��JWy���r)S'M��fO�Mx):m�?��*�ӳ��L�Q��j��M�~�H����Z�1�."@�����OZc�z�:ur%�@�HՉV����K�����3��)���X�_VˋN�JE�\/���w��1�_���eM<�箵Do�
}��_���M�>+L�t(��}��'�ʨ,!�\5�N��ĥl�閻�]
3*���4p�� ?�����i��F$��%�J���A�)-��x!2x��vt�r�V]]*BS��� {5���{`>���[�����AɌ�I:+ډ���D,�6q��bx� U����l�+�Lx]1�F^ţL�&�Z*UF�H:��&�<J�H<�ݨr� ��T��nCݯ��+Z�m���<
"�	ۖߧ�� �<��樚w�V<�gʸg�~lc���n�=AZ�PX�ݩ��VIR� C�\.^��뼤H��D-G��o���
�PNϪ��
�@JW&K_ֿR�/����3[��׋TЋ����S�;G�ğ��&_Ud�Wゾ� z��n���=�G���x���ޏ�t4�n��

�[Kx�#�H���) ~����{m�!����nr�dv`�9�S�«fL�
�k3��o�G�qt�u	˴J�j ��9[B�.q=~W��S��T�T�TӇO{Ғ��B�b�/22R:	E����I���41ɫ9bP��q�����|m���0T�����G��a�ܪ��	�Co��`����:�2��v��/767M�ޡ���� c�-<@T@�D]]]:	���fO.������t�@0J���3�q�ۅz�5� ���LQ�4{T<���mc�g�WyJ��8������4c'�CH bO2s4���f7���XȗG�<�����][�;��	
�? f�3�OK��/�a��/�QJ{{{�=���ƈ�qNzM��_�TcJFFYTT�̟�=PƷ\#YQ@����]��v�>����&&&�T���dW;�oQ�uG���%I��)�l��< 1��͂@�0UTD�߆NO]�GFz��B)\���,�B�%2nb��XP�Yv�`F�D��q*AQ;[�R����UH�t��X6_�Л���NwB1�@+�0w1��&Ahꙛ1����Q��)����)c�v�ˮCA����v`&�W6�܉�$�)'^�����ܒ�T:	��4933���j���T+��xw�i7��I4UK����Rݨ^�/Ta�%Yg��>�뀥��Ol�:�$@�VԎ��/���)��Z)��Ajũs�[-ٔ�>���]���~Rյ�Q�{�Yiq���.���,�$�	9Sn��"�=�a"�B� �џ��M
cs��3�a�������Ϊ�vِ���f�?e����A�W7�l��ˍ�$��ocs�,�5����V�jz6ɰ�%ft�#�B�9��	0����4������l=W���ͅ�X�	f �8���t�?b�.d6]��߽w#۩�sz!Pi��,U}�(�����>[�# 9��=��F�L��fd}��F�}�!F�g����Y���5�[��}?�
��=\��չ D	��̳4�ET������G�'��G���&�:8r�����%��5�;��
�Hf�����c'nTi�Ǎ�����=}Km�g���4���!+�a�m�,����������ڝ�݊�.R�.l�p���}PwQ�6]�Z(sR��t�o^������B�]�h��-�G�Ӿ��ck�nުT4�8��f8���)���V5��э��3�	+�'v> �&8���?F�Ds`3D&W����eZ�>b����6+��<��ِ�|�Ʌܘ�f
�LY#q�u	/���c������m��&''��<�}lDs��IA�/dc)Y�o]�D�[�o6�����ON6)�oL�EnVӮ�0HҦj�}��#6�����-6q���#� �����PzU�$w](={ǣS�ot�¿��06c*�a�2�G�Ϸ�(����J����P���3�ﯤ�@ Y�M[�h�.�B���ƀVk>��0JdF߃A�x �ݹ��E]W�o�F3�0���⌇j�әCJ(�ܟ �0�j�'�Bp<bG�k�U�H���c2*�Xs�W�Nx�}�x:�*Xޜ�I'u�����P=�����AҲ�@+���#W-Eq*�$#?00	Qa��y~oǓ.�'p��P�X@�L��Uy%Lፇ.h��>���[��U�o�'5��B�bb�fgu�f�+���88L����۱-p�z�!���E�(���X75�' �C}�#��
8:�/J#��H�@��)kNN5�"��6�ss��^�|�H�x��|�U�#��Pt�i(��p����e���,�u���	%h�
���^���;?��	�� .�\F�"�B$�� *�;�M������l�ȯ�Xf�U�H?�q����G_���3��M�~�)�퍒�2�2=u6��Cc�*���)�h�b�a漠q1{|\�$W+zn�&)��x�y��Z�$#+�9�ǔ5"V$�yqwP!�~rԎ�d�?\��w����Y��>�����	w��~x'���M�j��wL����Ӏ��P~l�p3��)��눿} I��c����P�Sh��޿���6`%0O"`� Ǎ@�,Ć�p�p u��Sex��P�
��>���g�$�4���yT��Օ�O�����Fr�d(_�t���\�ȕ��+J����Ų���Ñ���{�ր��_�t�����-��Xހ�b�:|/`*��o�������n��'�N�
�c�����Z�;����Z�8zy�'���B�`i�G�$�i �ph�?�x{��G[8��H ��Z��ؖL���aYtD���P����A�}�{���p|����b ���|��<4����t�x�ѽ��{+�	�<L5��!�W�}Cd���b:�p1೹k���g�X� �{\B��]%t�2�'\���>���:�'�B���}/ ?����`�p=�H1�N9��h��܆Z/�J�/Jh�����V�؀nm����Ø�w�ޥ���8������@�q<{�����!"b L3�4$@�;skn�Zl��UYU�9��Ks@Δ��jrA�"�նv������Í�Z���j�,A����QM�U���<V���}S'-������r��:���:�|FnO���B�Ր���~cw(����	�E�D_0�\p5IUӗ�HĪ#�iGu�,�ˆ�˗}|����T��gݟp@����K����*�j��k�ɮkb�G�Շf\�ԗ������G��||f�'k
�[ g�y倮"+��Jv76F��J��8�e��T!cqqq9]���7����9mfx����iE��%%��/��������Z�e��x��{���$����mEꅫ.Y7��1W�I-t�{���i��<�[0��~MCs�p�C%f�(}���Pΰ�(5���D�RR�c�5=�ש�ot:� �3�^g� �w�[7��N���tP����\ŀ�����F�q��˓x�T.����@dxX
�0Yt_st���j[�$\\�~��lu�H�ca��嚚��_�,�ѽ� �T�A�S�҄NN�ņh_A��.��Q���%��NΞ�y����X\�-W�rJ�&\�F����;��A�!�Z�w���FzU�Ѷ�oZE���NW<8�h�5���@�Q5��.Od�ӳ�o��|���x�r#�fLƌ� v�V����:�����&���ɻ��N�z�������_-Z5@���b'��-'���/)`J�/���D����^$α�}�ȪZ��__igL=3��f�c��(�����v�D�0��ҁu��}���rƑ��[X�`*�;ġ�6�X��k���r���*�V}t���^t|V�3777p"0��V�c�Q�k'��)��:g;h>`za�����ǔp?>�� �hih��=�ճ����'�.�a)�L�F����	���4�ޕi�����~pu���'(6��]E0qP�qB�3���hc�4^'���-d۷4�h��ɺٹ<^�k�yn)��VQn-�]���yk�x,�dc��<��"$"�&�xK�x)�e���/�1cb#
�Ca7s���A` c"����uY(����,�4i�*�뭸�x�ƌRE�9,���
��WЉ���t������]<u�|7c�lA��w:�����Ɩb��W��L������׈����B�g/�!�Ev~�t�������s�m.Cn�]�p�ͺ �}S��Z���ϸhl4��q�nD�����U�9��f����B�.xd5
�S-S5�9z/�_�7��3�#NV�!�����GB�T����������kGNg�%y���u1���K�BM|�N�\m;c��G�ط���.w��
�\�;��d��y�;*�Ǒ�)4���ƾ�^%��e�uN������?�,1�#��k~e?�޲��"2,�k\~/E��
W?݈	�f�����i:ק6m����c������͢oV��M_֙Y���Ӊ&�ş��:z@��.�6�z^a�'��gzl�|���Uԫ+��h�<&�d�w�-ܼ-��va�<@9⻹)zZ�����C�EޢY͛��Qw-�Y�HwL�mx7�ל�iY��Hh��ն1. `k:�?��1�k߽�i��ۺG�LR�ݵ���i�zb�s[�O�tzt��&V@TɊB:����j���l�{W�&�$l��2-�K�ܧ��4<^ԁ3�����X:I��1Z���
J'����}m�t����"rf��zV���k�Ǣ�k�wS$O n�;��������'@ٮ���.�J	���my���j����e����P�5�*Q���hV���(�d,����`no�&´/~^�>|�o���"�:�`�~ӲRM�c��|�u�Sf����t(��h�ݐ*�ȫ����a����!�q�!v���s����n��r����o
!t��H�@��9I����~��aM�<NK���y���o�h_1�����	�f:����
j���=��w�G�T^ڻ�˺��d]W_7��c.C��C/�;~��r�O@ӈ߃\^�%aj�,`�2���i+�;�~W,d�����[u9�ժ��L�!Jw�EԦ��&z��{&T��LN�*�z��uW�
��/!{������<Nl�cp�|_ޜw���f�u8�����w��>H��W�Q�%�oc��-�n��b�Zh��ڭkkm�ѲBq>�GS>�	�_~�/ �ݥ��	~�,wqq���B ��Ę�O�~���T�6+�Z��*��w����gK�(����(��!-�.�)���D�|5�)@�3�]Z��!�Ͷ�]����8�_�N�/8���'T�������M%t�j.�x�K ��.�g׶�l,e�G�j�`���yD��Q޴���;����}�]�(�ܙ�n������\:*))I5sE'37s87Y/h�����<e�V�o;�;�2"������B���V>U*��>�	 �mG�RR=(��8��
�V^ˍd��)ozIy����̘�u�y=v�x�Yc2�R�9�4�� ���}�Zg8:�5*�N%PI� �\P��M���Œ����'�(���"m#_7}�����7+�z������������y���*b�W�n�xNK�ET�_�m�{��VT�U�!1j$�U�?�϶����1�7K�X;͙%��%"vp�bc��f���v��[NF/�g�)�c�8��ʭ�{��!;.�b�V�}�"ވ��T�H�ڴ��l722�h���Qk1�Gh�#E���ʘE���_�,~#umQի{����Ô�D�zBH$�`է�1�ᴲ1=�')r�t�-�e��P�*@�̶�z�zX��5��x,:�.�v��S���<:u9=�;��;�{W1����xd]չl����jg��F({�;>,r~���ț���H��H�̴L4c�^ Wӑth�R>�S�Hz8H�1�6���cQ>Ţ�P�;�����d���h�r�)���suuu`�k@Kp	���RŢS�����lo3��(�'T�Ƶ���{�|o> ��My1���:����'#UV��$$�^�~�R%S�d�H)J�Ȉ�����:���=�n9���WְH�F����VN��!v|��,�� ��7=L���5uĜ�4��V	Ԗ��Ą����g�V���t�zw��'��~]j��_�-#����|(�(G.�'.GBF�@x��YH� 8��  �a���v����o�O�S�{Dw��~L=�@�:A�f@y��B_ӌ�ׄ�"��|ˊ����ί�c`v�e�����~���e�:�ug�b��}�v��@���H�A5x�H�O�������ɴ �p5Ɯ�}_k����D���(�`ut@�w�g|9Y3�k�۪l�����Dћl~�e�iS�U�x;�l�	 ���2�>Ûp�s*a�6�� /�<���N� �@"w����X��s̒��+�%��_���Wqe)|��Q��
��F�"1� Q�v`�vW�;��"�0�!�}c�h�C�k��=uY��"l��w��]�n�h�d��k,>����P�b��'��:*ʮ}DQ��0H��nP�i���TI��n�T$j�a�����w_����?�Z�Z���ϵX׵�}�3�c�=�.�5��vTA�YE�w�'>�oK<@L��ۻ2<p*�k������#i��>��@��p>��a�e����)-��-�hs�e�NFUǉ�J/>Jb�X�����m� ���矯O��L�6��R�l�
s2�zc
S2���~,�~�w�N�=8��1>L<��i#�fF�Gs����7���f��}��g��=|�QUQ-#Z!�P����E��{&�������N�G
	?1���H�@�5�,��ZQ����Ѡ���(�:SC�k��j$�\�����9��)�[�<� ����� ,������#��[v����d�k���`-�;Z�?�N��c�V��mb-)�����o�|�(4�(&O�?Q����s�[�6Fg��Vr�[��C/�aZ�smۯ���HWM��s�7��������N��9R��])����`����ɋx�ߍs2 v�A}�#��ۥiq�JGD�c���{�$�3ְ,�����㝬�[�� �H���x����e�c���0�v���q�����Ց��4���|(;���`
�$����ߋ(�0�Xƙ�85-E� tb'>*����?�֩&��n�Q�	I�k%tLG���+1�B1��qDQ�1��	��`�b��A�5 �@��q�뙋2�Up�o�g�4�V,��	�zw�}�%�}�l�lxs�M��kn �Pl�o���Ұ�7����ۙ�_r��;h�~
bD����. �XI�.$�B���iՄg"e�I��H��T5.�.]9D��e蠸 �,ji^�U*2�=�|-G#A�o��S��<Ya�����҄���N�{"S+��@�R��b�2��-c0��ޞ�;\M�W�lL�+ְ����v4/s�3&UѸ��W���9��UN��FMs@��/�4���ݦ:@ݚ��@�ħm�������6gE�@6�����������IA>&�>���kaʎ3{�-xBC��<$��qf� m����T�-C�۲C������|��^50�v�hA����_����-Ƭ���Mm�&���xF�ã�o-���&\�ui��~�_+_ 2����cH�C��ޏ��Eui�q�*�}J�H`��Y�5fB�x�i�A�k+@��"z5��2��
U���)�z�/���P��*�@O���(��vf����+hˬs~������NBbv/k��}9��I-�:�Q�� b��&�G�-uZVM��	�������4S��	(�!�l4Sϵ[�m�I=�S�����?��
�U�6�[|�˔���^A_K�Zoi��i�^��xkN:�Fb���7	j�a�R��*<^�*S͋�/�:�0����X����vȎ�i�R��#���ipL�y���O��&@��W�Leqׂ+D��ZMXO��4�>�����j�tdq���eDߺ��4���ʖ�7*WNʳ��S��>^���G,��������3>�(�wF�l�b����1�,�$L��ȟ �L�`mW����]���i�9�!vT�,@��d���ŢM��"��Q���Z$�q��|��W>^.�(K��Z��?Eh�h��K݃<4�Q�^��0�:b!A����N&��M�f='3�wV�qhh虘�C4^��
,/�gE�tu#߄�_�`V���%Y�c_��SϮ�h��="��퉻*~u�E?��#{d֌Ú��?�tb{��K[CօxA�9�"���)Ez!�"������_��D���A�J]������Ev��-t���w��iH�\ӧ�^���v���{X7W�ρ�\�:�;�����pvj��o�x��8�=~_�Qm�&�����l�O�9�t�s�˪�ۗ�%�kD/����0�� 콯�z���M-��{�\�kV_k�FG�Ц����8^����uA��Y���77��m~Ԋ����a�/��0�H�&���7�<)�ìYv�
�d�밡VVK�u�;�u:M�wxdj�V�	�ȵ��u��0~*�~�q{�V��ap�W?��AB��T!�/N���R������������ϴ�Q����)�4\J�ABS'��?[W����g�ҋ�x��k/�'&������k��ξέӋ�I��NO'�Q�/�<3v
r��c�w�K.a�~�"������$�|J��DR[Sc�u
��m{-z��׮2�� U��C)�W\�o��~�	�ě|.�8{��Y��֯���fhΰ�f��$"uq	��]�#G���˓�e��gr>���v8�z����!��%�{��mu?��W��<L���Ƭ=�/*�䫪[mJRI��Oe?�l��٘1��]�C&-������a^'c(i)�,ef	�Q���:<�-r~��yZ�~���H�T(��s�C��I�#`�Z�`�@�ܭ��偁��{���w��۽�p0�L�#V�&��RƘj��3�1M��݆Me ��>�;)ٵ�:p��CN��϶�D��eO��\�^ �5�;	#;O�6gLcD��p�y�[��'�m�.�������^�!��������{cʴ��%�߇��|����r~��[���b��;y����#ޮ7�o�i��N0�$�\�3�����kQ~^���F+�:��f���S�cP��Eb�,v��Q$C����$ʞ�+�3�fo����[+�����.�(�A�I&�Ȓ��uj��QSC�DӴ�B��$�q0��-�'�,��~�&���T���rg�_�H�(���B��"sv4�0���y��_����Ӗ�ym�Y�
�Sf�SK���.����^V��'�+��viniF\8��-	;�Y������qEb�^&`�[po��K�^?;*x���5���߸������ k�k
�+/s��k���ՙ��'.�$w/1OA\��g��G�2Sw6�X����x�~c!�]�[u��mМ���?"�}�o�8�u-�t���#9����ǳ��/�<�����N��)�3�@�Ε@o��]��� �$�J����&o��X���<��Ua�	g������V&oc���g�N��y2Xn��T~��+�i�W]���(^1;_"��!V{�'8�"��ߔԒ�9x�k6o;/�L�M&��3�8�OEX�S�ӀI|�{����y4�I	���V��0<�r��F�u�j��q&����G���7�z=��!
@%`J>��	�&?��/�o(�U�Xv��4��U��FX�ȭgVS~���X������ړc� ����y���hqS��~խ4��?�c�]�����3�/19}��Tߥ�/�F�/��j�d�zθ6�sI��� �1J�p�"5G��Hɟ�|-�\��1i�t�Εs���?���Ա�1�̤�d����׾��:��b]�6���|���@th�j�|u����i�ω��2}�b����i5NhS'���G����Ľ�r�����y���iG���J�dyx��g;"�8oO�{�ߕڙ��cL�_~r;|�.^fֳoI4>�8��sJ��D�f��Ay˟Le��e�:7K����Svꙅ6����G��'sV'�8�I��'L碵'&��x岕��ʹ����/=���ѻ{�򘆛]�⁠Ԍނ����׿�.PS���,�ZMrJ�"I���ygq*e�t�Ξ�1�(�V�VK5��U��������Y�a	�`Ɨ�$`mV��2{#a�u����5�.+@�V~j���3�%�͜��S��?m��U*�	eƷ���৸���a�v������W������R��RO"Ak�C�}���[�5�s36�'�w<��	Y�_�#%.ua��$��Q�ы�o�!�̗nl���ߝh3��FGS��iXpǉ/�Z����tsv?�8k�;�+#Vj���:G���:YI�YؿIe���Q2bI�ӥ���B�v�uXO���E��������;,���nC��%;�JՅdA�T1�����	��pA��AhKa���P�������6���L�%�����%l��D�nڤ���T�X�,��,tx��x
��ܷZ�M���́��C�)�2�����B^�|�o��̀&�M��D���:m�����(��
����z��OCg����m	Y�KB�������Bw]P���MlRwSPV�T�}h����Ƃ���p� ����9�~O�_��mz�du�@���i����S�ى�K�f@����8�E݆>�r�Q�����+O��?�SRS5/���S䑩'��q)]L���k��{#O%���4�����X�c+�`XSrZv�B+԰��6�ia��'�6���V�+��Gz�	p�TZ�lAo	���mc�n���>�u��x��N�7N��	�凜�03?]���������c�Yv'� ���`�O��'��}ۧ�z7�D�<����`ƶr���NN.� �?��i��}�2X+0	ET�����i���d0�N��|�z>B�@�<+�� >ʅ�w\-�9�F�9.�B���Q����H'�h�
G�i�B�mG�Õ�L{J&Ŝ�}��a�Ё,���n����7�zյr}@���nY-�h���u�Z�<]s��_�ࣂ �ţ:������aۻ�u���m7�LU�ǝ�XG-�Е�NȽ��>�Uom�ή+�@��W,�z
-C	}�"O�'����؀	5R�gd���ni�m3����7�����w�7lE��(Z���;��"��j���"�C�Ⱥ&G �Y��T$�t�sU�cO����S�׀���w��jv�u�ݥ��\b���r5?7����b�����/3v@F���}�̸G? M��A%�d������̏-!���{/զ�/�`�Ґ�Mَ��D@r�Wȟ�b�w�C�p� �z��5���C �:Q7��젼U�N��6�4�J��į��z�~	�5�%W�	��J������y�Y�T��&�� �Оd'H������~Tq�h�0��/w�A�J���(�`!�?��6�(������X�A\���Ο	�?`���@�jޮ��=������?����y�D�R�<Jw�X{�4*�����^$��V�n�jb�W�#ޣq\#��[��]�:$��a��V7_�ox�1v״:�+�� �}w]ɾ%����XpA��w�ݔ ��y����i%`_ޮ>�T��g><�m`fB[��M:�2�U���c�L���B=3(�B`�7�o�]���44��d*����TW���ǏWu����mm�gΜ)��|8??��ãca�^��,����]Y��
C�a�Xp�9/�Q;����DL�3�� 
7�L�o_�\ �1.����Ұ�g�15����r�˗/�YXJ�ƞ�+(p��ܸq���J�ٹ�͛7�W��t������r��ƵϪ��PRRƤ��MM�c����7�t�0�iN\�l���n�qr�z^QQѺO�e�|���¢��$)>>5�.����e����.�=�r$h�*��Qe�[I����3����-��5"�ovޝid0�}�H{fB��
,�app�v�x���)*J���9�����x�)#p�,���힓���Ņ�B�Ar,�����Mv�{�	9��T��u�*���B6C�U]�򪫵�})�E%%-�;������;%��������|��r��U	
�6�g.�,����L?B�0;�g��|�9f��\�cq@�a���5c�&8���q��W��E�x.'�ZSK+69����W,2�S�1��Z�5�J�&�����jluV�f��.]ʌ�1,��k�'���㶗�>��_��cm5���2%�ѥ��%sYs�� ���B1*V\�8R蜃������%X/��ɕ�JfP����~=}y���4,�������R�Lpk��_��z,�Í�0y9[���������h�S³�o|h��rZ���q�ΈL��&B�?�DU�����ޝ>s�lQy���B�}��0�;u�z��[�q�F/=�g�b���4�%�Z��|�./\�z�W���DY���|��R�c�QWS�l�r���o�����W!��B�z���NSP�`:C?}��Bl&�����%�X���u��m3pw�[}�#l����5���v��w����S�-p�c2�G'[I�C(��/3SMI�<ΰۜ�������#�'�iov��#`��P��I����#��� �彤��W�6��/�?w{�%�^�c�ۥ�M� ۂ�D\�-���;������RTQ��(�X7�׳��P��R��5�ORFD�*z6b���+a��Ф�P�s����X���de;�:�<mU�����zUwm��s����)lYܫ-exDKY�W�B�/w��@2MW-��\����#��'�bO=,��s��]��㡦�]Rޤ��f�K��\������)�!�I0�q3X^���mĤX��n���2^Ƙ'��Rx���R�G��m������0��H�o�dJ��^�xE����p��_�$����R^n�X�>�b�x�qY�d���Zv���= <b@{��hV����
�
ڑ�n�r�-���ˇ/��]�?���z
6�LK�J���yR���=7e&�X����!�� �N���a �� .�2SE�����&�=�O�V�j�������m'��ˊH�~X@���L��S�^�u�MF<��\�+|wQ���1���K55o��*������J�N��r�/����
r,볥�;�� ���k7*:<C͹�D�k�e���X��D�d3�͊\":�;�j�>I�':��\ ��s ���9}T-�����j�So�{ ?qw^Pl^P��{f06�{i��٬n�c���9}��K�x =˥U��t)������'�y�,	����rѲMX�է��;HX��A	6�����?��Yu��}��²K�gk~�O�f�X2p�M�N�x�&"�� K��Z }����V��o��	EZ�^T�Y��QQ2V�xM��h��$�a�n�{e�S�q��0^ch�&�C�r�|��T�NZ!�}5c&����R���g�Gی�<�_��h�>c�H6;�\ݯ�'�U4�`��4h�2u��'�v@%�N幨\N�&�� �kU.��݂<oK�ͦ�E�p�=�6I� eK��M�暈ν�����1���Ujr{I6�v,��"�S�#�j��@\��s�tVs@��U9�b��ҋ�Lӈai��H�0�{w�*���{�Gc�:��V��7��p��ޣ�o��EJy���I�s	��}+��(�8��5PaQWZ�Q��&"_U���<<л��ޒ$:�oAc�2��G�1�dm�/<�?0�7��u0�U���ui5b
v��l�m�hg�[l�ppܗ�T�=I���k�m_2�t�`��	h�t+�wr4(򅼤��X7X�5��Co�/�׮_&zf0��<����KN*�H��BQ_~��-/a�����Q1o�Q~�\S�B���H�kψG��cvt
���݀�"y��6�G׫0m�q_Gm�~|����/A��@������Z������;����d��2���vX���3���g�Hi1��.`����}X�(�T�z�F��څpp}x�4ʲ�5�޽�JA�kj����4��
 F4.jX'�NIsNWN���߰aϦ� ǷYr ���%�fn����]IC֟��Pu�)�ef%��C3��A[&9�4{�I�? ��0����U�{����G�>�?$�[���m<��eAM&�����b4�4AH�d#��U��T}Bxi�����!/���m����0ɖ�@�ݦ]��xf���3"�]��������ǰ�	3@�w<��}�v~��3�c�y�[]S#3��鐌��#h���	_Sl�S
UVU�P�j�S��T�G�M3ߒ��V���|�R��v�m��Po�y��|a��8p�hWU6s�#3�`p�mI�� �T=+���V��^㩇��D�l�Ǐf�Y'A�2m%I��+�]Y��l�����eWK�(/Rk?�94�)//�����U*�1|�m�ܲ�?V��غT��`�rK�xtV�tOnas���Aq��naq�2�E��2-F>��F��G?��HP9�|�����-_�E��sG!��{྄j��z�͙��-���t�u��Wѭ��=�QC�tH\%�{ml�C�
G�tp�ϨΖ�'�ʸ��)n�+p+��]���`�y^Z���F?�߂{l�,x��H������� ��@˭]7��&�������$E�ׂ�r'����ge�G�l\n16kk��E�I۠,�7�$�� �T�<��	I�(�V'�,���B�̰����T��� �������ws#�]l#��?���zm#�bM;����/p,B���q���Y���'}�Ov�_��a�c���E,�M{��b6�Hw�>�,��T<�A��ON��BCߩ�ORwm�����=��$�:��x٦HO��]^1M�@�-2���$dW5����wkt�������&1?�>�%	� �~-䚥�)��%I�<�df;g#�n�xWj���Κe���O�_lh��ױ�K��6�W��6_f�/�{/3�z��Ӝ�mj���-�`Wy�.���PX[�2'|�u��ʟ���A^@K���j@����/���2U�MR8���b�S`H���	�*��d6�W\WC?c�J�����3g��8RV��M��}������}���x_�՜T�B�Wn�ъ�~O�y��Z�����&�+��5<��:������h¯H��7�}��o�7�i� &�E�� ��gsPE�I��i-����~�������QE}r��v2�:��Y��e|`�P���M��1��Zby��٪�ißV��|>G��l	אg���-�ɝ���Q���e[P�K��7f��:B ��T����f0��������z��m����׶�/���щ�)����ֽ����ۭ^u�"����/���4��жڰ&(^9��J���p��-'�98v���j�;~g�R�?����s����g�O��|s�J��ɮ*�N3�}�9�* q��9����B�-r��-���tr���c�g�:�t��%l��SGE����$���������8�hw�c�$�7�y�4F̭K����3�C�Q��l�������h�����<NM'�Q:�������?$�I�F���}c!k#}�s?Yw��~��3'z�`�0J�'�eOD��NA���ΰ������'2fnB�,�<�����l=��Շ�F=i%-�b�U��?��OV3#��?���[��ēW��<�ժ�J�_|nkR��6�%,u+o�������م�[������?B�G����'��<t�ڰ� ��OR�p��0w�S�d�4��>�/|2 �1�\3E��K:�I�/7m.�+C@����t����?b�|uw+ ��;|�V����7�`�&%0�\�dY���p�U����F�K�ýw
S%� �P}�Z�Z475�Rslk��( �H�(��x�˲J�@<'RsU�є髈�Χ?ے͞���c"��K�U��%��{�lYǛ��y��U�@����i}n_Zw1H߭X�&�KY�Ԑ��s�W$�>�Jڦ�}��T�c�+le�2��]�qU����}���K��>REB�G������Z�_X����+�l 0��3���	G�:������Tg�Ro`C���oV!��+ k��}���f���JZJ=�Z��z w��e�����1��mr�eƫ�A�Y�F}.�)ˢEY�Vl"���R��#���L�};��K���K�zm�Z�xtx<�x<=��� ;��u ڎ=H�I=�{�8�Do-�8������%�wrjt������{$�8��C�Z��-2=eBľ���������O	2`�T[�?�L���G�6�%�,^���X=����"IG4��M/����HF���7�9�y���t�
�.�5�ODW((TF&����>8x�;������DU���"@�$��c��߮%5��r�пv��P 9�'��?Ñf\W��lq�� �P�{�G8N�F�d���M�.�����cHA�Q�9�C�,s�5�M)n��d|�ғ��Ժ�CUd��c��֫�g<b���v�����uK�$�ZzW�}���;�	r�5K.[��D�/_������ݟ�=�@_�u�"�k�m�%�d=�˚�ЊOrwC&	e�|6���h����	�Z���]����˧��ޭ�p����e���9�TI��濞�[zI��+��YVK�&u#��C!�/��c��3�f��TN�,r��h$d��z��'Y�֮����K�;�;i:~�hT��S|��c���b���j��5?h�#���5��Z��qmv�8ȭ��{j����~�~�6�;�zt�0�8�.��b������`�]w]�;S(,���l;g��F��-�Lv֎��g���jHS�=[��8-�U��¢z�����Vtsy��� ����ρ;��TN�b���+�ti�}���nM�e�^T*ŉF��U�ʒJVm&���Ms���ԡ������񑞿{���Q�@�zԁ���$����N�{Ē��IemZC�����U�i�߽��yH�˖Q���On�=���=Bqw��6���_�E���_��-	0\�g����s�~�ZeY���i����i��U&��j��ޒG@��{I�yM�1��xw��f��_���k�`Wǁ(&/��H@6�9�$�����9Yz�)�aS^Rإ�tT�u���e A����#aPY���z��vu@'�v�Y]z	,9�U���`1/'���._y���t��U;��HV@,Z�X&&��6����Vb�^OwVY�Q�@���j����ة��r_��.��!��?[w��J:.>��[����1��	w,���(�Ue��
�"��y�ｙd��Pb��2���b����K�M�KA�9�%ȯ�Ye&��+
�>=�UNU-#}g�/ӻ��:��u6a�Z������^�����	��t֩�e����L	�CA��'}��w֚���5]%��O��"@�B+��7����VbV�VdT$���n�f�|�on�4�'ō�}�F����\A�βc����驓���� �BǿXtswB���S]�2T�	,6������@ɭ,d�������ĨeB)�;.�f2��.Z�5�����i���-p ��vF��U߳������E���`q/?�����)]ޒ��j�X����߹2��VǢ�
Z�$!x��j�WT�;��-Mz��7B[��,"��U��]�����ý� �+�O��Ȧ����\Tk��?�Q4>���SI�B���W�-�{�M�)t����Q�Wc~	8������=�+�\I$%�pbA�H���]�&�w�[L�Hx���D����
�,�й�q�Q qDA@�_���ѣ%�� 	\`]��$@A�7�
��|sLzK�Y5-!O������%���D<b���c�8�d��ײ��'Y��w��R"�12�az͋�n�E�8E���N�?V�Vgǥn|��<�sAM�Q�k�+�P�H(��������n�	l/fr�b͞�C���D��
��%���+.���S�l����Z�A[�B.�����)zK��>G��d��L<q_�8�n06j�~V?͘�r��R�a�Kc����5��{$�:m]��k*Q��7?�x���e�]ݰ��ձ�d���;�A\�wρE"�[F?���C�"��A{�ի�Y~�g�4�3�_�ԣ~���͡ֻ<�F�A;����D�у�3��3*��;Y�1�<��D�V���l���0 ��q�د�[�X�ļ�n�q����79�d�O�h]8n�	�<���lUuI�n�nE�I�$�/�X�N�>�ؗE.�w�sE�,!En��~^YDl�xm��cb���O�RTWt��w��(m6nml���|r||=E�A]_˟�ci�j{���xo!��w4�x�:�|�I��Ol��΋D����"��j���ȋ?����-�ad�rX�8��uuz��:iW�Tk�����_b����,����*8����ﷅ�˳�~)tW쥚u��|���-��B�iw���YR�H/�H�cF���v��M�0���{|�_)���/#M�ʰ2�S5Y��
�i�Xiz�Iĭ�Ѡ�#��K��?��y��7�9T��NRQ�����m���RO)D�
�:Ղo�klBK�<R�������F����d�q��~z���h���2*���,y���U ޑ�����)�@=y"����"YM���;_�-S�����8���*�)�z�+�HDB2�G=K�5G�w:��ԯgX`�,Kc��|���eK�rqZ�^n��B�7l}o�V`����CҠL��G�J� E����dj�eޘm�o�u���u���i���>�a�N`C+hr�����ȸ���6����o�Ĉu�$|���X�v��Ħ���\^�Dn�z�T�)�];mwhcU�X:�a�*�Qr��i�8��>A�`p(X��*:
�qZ}Y�yqcK���� ����Dx�"�1��o$�k�@H����y^=�*�o<��C�� H��cًrY�k��E&b$^�m��ۇ5e��@/�O��r��ɖ��
�����j
�������	݋�J�ψO'����������J}s�l�R!͹ض��L~7��;QG�&xO�C?�0I�K.Hb	�̴H��V�$s֨�����d�?�o%V{�d�6�34��oxek� :s�p�,�Gh�O�Z=��i�Pl:K�����AQu�Vjl�� k׹���:�A ���/�W��1��}��`�K����b��V.��$����6�C���<�ڂ�P��{WU��~�Ay��1X�o���Ԩ����TK4҂v�恿+�4���U_���"�p2b��`���3��I�P�5�KKC���KsN	⠴\�t^'��<���J������΢EcL�#Hl[�!qcq�K���2�K�K��F'o��Rw�T	��QEn����yQ�dhm���J���{�k�Z�qѱE��5�H�=f{<�4�7Xϋ����L���v%Fυ�DU.^�%�Ԏk�ZA��H9$!҂)�f>~�E��c�Y��K{���Q��|d��K�D�U�A� i�����ҐI'?(�} �v4�/*Mj�g���.���M�+�Qyh'w�\U�J��C���,{ﺔ�ӥ��"I�[�WX�翩<U���[u���Ӌ�����:��,ϳ�*�l�I �Y�+Emw����j�f�FP5��Խ�Ƨ�!wyR�l��E��&�.7b��k��Y_)��^�>0����������YP3��V)0bV���/j�K�I�ZiS��g[��}y����2~T�,V�JƁ��wZ�*�Xy��}@���t��(��i����� q��j�c�IE�Ų ��%ع��������˼��PI�+t R� �	rlE���C}EVWGJ�j���U~�OOϼ�XN�p�٣���4��(�]��f�?����{��8���̏W�j��� �-[��x�f�Uӹc�V]@`�%wZ����Rі�vj%V���۳�>N7��ݵ%&����쎒���]��5R����zP}b������;ex�f=�D�Ŏ�������i\vT�J�V
rG��v_����w�H��{J���l��a�k��䜏2n��Ë���zaX;ꮔ�!_?��b`��Rb٧Bl/Z��j;�n�����hjZ��J�Q�h�$���:�#D"o��j�>���j���ρ����6��{��/��q�l����V�l�)��
=:��-��g5)!=�pYvRyy�>I�+Q���E�N̋�?炦{�6sO\yg{=O*p�)S�VVJd�g�d�E�Q�|hu���^`�Jq�PF�SQ�e�q��=Hn��ǽ����&���Z��=��޵�7�)�<��Kp]�;�iR�8�L��<`�>�˥U�H�Ұ�a�k0	Rn�&U99EJ�n�gZ�!��F������(��>�ڱ��7z����1�3�<��]@��9����K��R+k���\L-����>����oCD�> ��ᇟl6�����WR-p~#vm�����������,�0�BFC���������%��'�N;}��_M�(v#�]�ۛ��T��"�1E6Y�W@v#JQ��_�C[R�qb�Uꤘ�'\��}��M@^����z���M�/��8w��k|ӥ�a�M���%��%7���H��͟��zu�� Yװ���#޿���ɝ=���+R �Q�zl�=�M&F���W�|;�V�����[	�~��޵�k�ͩ&��.�M���3o��e�k�vjվ��.�7�#��Pذ~\أ5S��իO��tS���5�C��]>\����{ �LH2P��d'&��)�F���מQTk���'�����w�ayF�uQ|��H��X��"�ޯk5�m;�u���|�~(Rdq���6�%�t�P��W.ۘ"��o�e�g�r9o�~�T��woޢ�ㄞ�$W��)^ _Er�,@Y>&��f�S�C�*�6�ql�k.�"=�0��\��n��0��A�u�'�K\:�c�uoPv���*շ��jk��x��i����6u��r��z�X�������]����4����H��y��mI��N�;ȟ��dr��[%0��/���Ɔvut2�q���p_�Rԅa � �g���w7�ˊ����<�-Kh�Ӭe�Nm�8��x����gF�,�Y�O�{-]�dbK�ԲF�����4�`6*G�1L�p�6�T�p���w��c����`��W�*�T�N�B H$L���C��)[G��\�����t����H���H:�v��K��6�o/y�M�b�R'�
����*Œo���!;2�{�ͤ���՟aY+�{蝌��m�|���+֧ʞf=���i!*�E��ljhvhc�u��[�P@��z��ΧV�U��;6}����u�O�UN�����e�(sE�54���\nI�f��#/~�f����^Ƽ�w��$�s������3N��`1+hꪠ����܈�+N�"��#���K.���TbAG�[�}Z.��bZ���RV{M��[��� ���-F���#�o�Q�!"����|l�؀� }i�\x|�A�*j�ƒU�ʎO�T�]V)�m2ަ���J�Eyٙ��K�FW�/k�l��R�ZQ�k�)u��c�[I���$e��J��^I�����_E��H��d�Ƥ����Ga+ MI���c�U��i���.�ϧ���V��)n$IO�dt݊cm\���Z��EE��&�M��	���C<�ip��4Ȕ @1�7���π�h�!<�$��-Υ�m�J�ߏcK/�J8��iTx�s�*6eW�kєQ#�ǀ��{SFK����4��L�A�}��9�b|j�'I����%Gl���n���}�s���ob�R�> 40~��&kh4��pr�r�+[k؄��~��k���'V�@��Ma����77��d��z�$IF��Dn���}�nV���L�Eh�[o�8E�n�  $=q�eR�;�wi1:��A5��3yO	!9���װ�p�����-|0�bS��k�K��m!�o%s�=��5��|�����;u�A�����\c����l��%."�A+(�d#�o볍p�g^�����^��8�&eV����73�79�Do��7��z���փ�܏��9�?����w��G�N�ש=�#�g���U��F|
�22���nu�p��G���R9R9Y�%O�H	��˼��C�fA�I��?o���T�߬4��juI��M�m1|���
�B�$ZHyX#*S�Wz��Y�ǌ�k�D�#�>SL*r|-��VZ�ek���n�8Cr�gMu-�q���bA���Z��)����j���v�����	�֊�+����u=�ǹ;��+8�@ޫ.%�����e;��{[�����1�g�~>�W��_P�M垶�o�j\vs�7J���c᳆p�q�^~_)�e���5�����Ì�^����w[>��1��V+?ل>w<�N�k���^���?:H	\{��'�cQm�@�7K鿬E��m����5��{�ߓ��ټ����46�[��'\��W}O�$`B6�wd��K������Lܵ:���jrհ�ص�3'������$����$��:,�b�G��J��XZ�6���]#�HU�Z�GO�PV��9�\{�A�å��qE�4)�2cf�����Pr��N�롯����9��
?3��c#B$(��H)w���'*�å�:���ӫ&��:����DZc�n�䭛&ց���L���WM?���f����YT���W��\���c��T�ܫ�@ �7�.�hr6��3�����#�ʯS1���{��]yd&3l>���EKm�ٴz9�E'����!`1������	���͸yy���z�i��qW4�}�Lw���� y���eUP�p#fT~�D۽5��mk�RE���wK9�V���w�}�B�N��?J�
��Z��JO�9���ޚr�i�)Ӯ��Eo�<�]8g���h�����S,��������S������F㕕�e�i�37�BK=��|��$��~�)�Sig|Ѥƫ����5��cy��8��������Ԓ�f��o�*����9/ֱ���;2���)��ٚ=�G5��}/��˄�ቿ�e${v�{F�z�Ȩ��$���\�qv=�Lj���F}��Z=�����k,q01V���xF䔨w�[�r��{SH�`.Z�"�]�7H�k4����b6}�,�{ʒZ�jL���]�]rU��iW��.�a\���TA�@r�ށ��:ta��A�'�Ľ��4�;���g�!Np�F;f�&R�^��Vi�̫�ϧ_��Mg�*�6U�FyC%Rn��bVK}z�?�}�{����E����El�$y ��z?�&,��}-5���^~�-O�DA��ŷ�jM��>��?��S_��q�X����ٷY#�L֝B������w{v�����z���m��pO��&�NEoKN��KT�B}�A���iw��i��|$(�!�m�4Z��6�h�;>���.\6i��6�`r��~.w��;�~#�V;_ŀ��\�q����;��)�T�<���*q�>-�ery'��������&5����WGE�}�
_E@D@I	ADZBB��R�v`�!U���FRJ��i@z��a��������޵��Ə�X�9g�s��g�g������I��/���o3>���i5�-� �M-��o1�H�Ӥ�i�387�#���h���y���1Zَε�`RfDgv�3�|n�Q�=���Uw̵X[W�+�UJ�ffg.��@a��U��*.��z'��
l��yb��GV�B�#�E�<��jbe%�\��c��L��u9�.�y�*`E?{�H��q�I�u���H7.c�1�O�A�/=�6��\��h��\ #�g�(A���5ў=�,�����E�O�U ���O�Ec�$��y���7V��i��6h���c�$/PH�΂r�J��!r�Q���r2L�u^?����B�����I	�k`�f��\�n�M�x-��P�\T�Ļ�L�G=tY[L�����68�6<������6}	/�/�<���W�V�?+��̵#9���a���'|��~DT�I��!>H��PƲ�@�ܳ!��ڒ�6�P��Q3��!�����dٹ���������%��Q�OF[;XLw?^/��p����YE���@]�(ϚZX�PQ]��Ǌ4��cD�J@E�"��W�8Ja�U��lz��i�Rq{�*��0p�B��-��X�6=^!�U��M��K��E-�o�j��qzI�?�8�vݝ!�������dB��X�)* 6�_S[�uݯ5�C�)�.�X/{��uf,b(�li`�����"Է�j��97\��+zh8��_��ܖ�V`s�u��x֯�m��WyD��kR�1�G����]b="Z��g�\؈~�6Ak:�a<�gR]�!�2��V@�;�Ř\��wӳ�S��ųq�� ���I��toX�3�e5��$5��mNUQ:_f�uM�c�6w�1�Mq$��3�U�Y�@v�~��?�����qj�����Y�	�ː!x���v�D�v���v�f/��B�>+��ϐZ9����Oٴkc}PF�&΢;.�oF��2k�q( ��[mL��=����|��*�<a���0��v�D��W�{�Ԩ@��;�n�9ܰ�AÏ��	ߧ��,�Ms�ݿOW���8I���{ ��t���ъ0�9S��F�d��q`(FS�*̙�<�H�'Z'��'��y��^�� ?�?[Ef�?��0]~1�-��Qqx��V�+��sˋ�e��2��͡&j�I�O��v�pcteq���9��(<���0v,b:��������4��^��iR�����/'![���i��(�|��O'q��3.����,ߋB^��n�䑠�u��ՙ�S߄�`�N3�O�1+B1's���c&���VLtW@�g@/�j��+ue HO�r��-J�*C��ÚU��Ȓ2��������-66�3�_kD^tQT,8مT0����֗�<k����5�/e���;�l=(#l����
_F�����������v�`W�W�;5��<�l�r7$��<f2�J�"��������Q��������ykM�A���])�M`�������Tt'Rz+��S�ZW��\=joX�������=܅R�~�I�N��:+k��Rf��Xy����k�L��Q����-W�\}
�C��-Z|0��os3ׁ��5���}��`��]V�iݪ�J�65���X W)��#9�В��d� P��a�����S0��=��<!:&����H8�y�Ə2j&Ԅסj��5��ç(��3��ypx9�����E�;|�0�ٵe�#���G;�ͳ����(�oZ����BkZ�����z1�m�NLN�x�r�֦�0��3��6/ߑQrGF� o�JmTL�ND��$s[`�X�*ێ��M_��K\��������F�f?�Gw�hK��y%�t!g�����,��l$�;:_!�d�h�ڝ���^\��4i��� 1�:��@�H��R��@���('�����[I����ϗ�D�m������ˋ�O��mq��\7����]s�@��rg>�.H9>���f4�@��&���!/S]�0֗���+�m����FgvW�kir����9s���C���f�I��I�id�>������T���8���L�ȼnf�Ԁ;b6,�K?6U��ae�}�y >����@&?N���(=X�TQS�`	�Z,Nu�� ���B7��Ɗ_m�t������GD��b5�vދ��v`��jnI�MB^�-�_A��I�%s���( @�p�C��:�����*-��8�] T�]�a�q��CK��ts��q���f.�*�#**|�-�P_8�4cኔ.^k�Kg��YkN�u���z	ږ��Y��K����/�g*?�N7Ǽ�CVI[���EPR{.�>I��oV���As-U��i�z��M��r��\���CkF��O/Xt��W�������b5>�
�S�,��W<�I'l���5�[7���>���)���ik��0�o��P7ۈ-�3���>�!b♷���u�Q��̰FUi��B-7�NX�*�eè�'JƧ�@���t]M.ҷ�4q�a19|/9��sD���hW��|�Q�޺����RŒ���G�A��G��̏�O좊��B�D�����&��bzP�8�A��şʾ���7��%����~����w�������@����&�t��b�=���vZ7�>�?<�X,w���<}��zt��J��?.��������!i��������#�(z��
���Ӫ#S�y�/h����}f�/���"�^j��mj��l"�f��D-x�G�^tU�gXǸ����"�_�:����ĳ71U�0����{�0g��^������r����徫�X�0��_���R�T�MW���5�yVsN(��9}yaǂ]C/<'`����m��˕��3�a�d�Y�]��)����O��@�a���Z��{�缡8��[�O�0">�L�N�D��T3��A�֚�Tn��5�I��"�\%�T6�Y@��+�Y�C-�"��������.Uo?�n���s��3���j�?�b(�-�q��&�5���ޘ��FXͶm��C�r��{����ꜼW�Q���O
�2�PB������|����s�3b�K�o���i&G�16Yk�e��,>ȑ�6*{�꤁0�ٽ��e����^@�B�>��ڇ䣀iv�P�g��"e�#?ؐ'���5�w<���gZ�hZ����`ҎޘHlE�������L����s4���"e���z�W��W�gѓr�Q�g�(�̧�=�HET8�زf#�Kpj���`��ј�������>�C�������a����-v(w�S���֝�	�����ΥN2�ϟF����,e���Q����M�y�(Ïm�8%.�G�O�}��(50������*�ӑ��쮹�]�tLًG��_�o`��r�%r�S?��v0��׮6(^�ۯk�E�7g�J6i�X\@�RֺP����,Ͱ,,Rk���r�����a/�Q,Ն�;G�tP9(5P��5�� ��xo��JY��;�;-Y|���N�3�X..T4�M��\�V$WD�X:���O���>�%�\�{{��
&�P}��;G'�wn]�1YG�U��U{p̗f|f�a��ہ�>�w@{f\p���p��{g����,�����cJ��`��)��$M�[���)s�kQ�sdI[nǏ�©FK޻�;!��EPNb�����x�{���/��D7��7�X��9	��Y����0|�4���`��y�S������ۮ6G�ܯ�Q������"�dA]�=l{�@]���e"����+d�@U�������v-�L�h۟��+��mZ:��;|V��b��y�?���';vTŏ�/�0XS�/3�;���.�ߦQ��d�V���4O��Z��i�MW�H9�U4hR;�ʫֱ�Y����U�	�}�]�Z��:4�0J���.���̇��43#׶��������� C�"�T ��e�̻�zғL77��uX�a�J�Z��W/��R5.#�?*7j��p�i�j_�b��Z�7g�g��=I��<"b����{s
x,^W�z��}绱,�;Wo���v|�iY��>}�@��	����4��dw���3�qV@���*��A�ٰ4��X�W��<��{aQ�n����Ͼ�nc�Ge��V�O��V�U��Mx��s�{s뫨O=�ɌȢ��E�ƾ�+֛�>����D�@=Y�5��F�]x��OJWU��W>�9��*�l�	��W�mIyLH��+Z ��/�թ���xVl�g���1�ͻ�CԩiCt5{����l,�-�$GS�,b��  ��n1�Gw��Y*����1Uj9���S�{rh{�{G�-���"�������	f:�!���!���������;����������m�<��i�F�SSC��B�a���0���1���cĜy�ӽ/�}���JX���B��ӣlh����Ej!O��G]�j��㖝�v��$���FK���h���,j`�y��JP���ww����"����BR#�ڵ�\��u.���q`���ˤF�
S�B���2q����wT���6��*\��C�.Zc"�}�_i����H6�&%î8uR^��eOl�?F(���G��ܢ�Mg!ﯞ/@�3h�K�й��R$� �Ǳݽ.�]xu���2/�᪱���e� qs�
�$M����E|!��)o�b`���=m�G�F_=��<ri���O�X�K���9ހd���c���1F.�!��u����@���6�1db�ߺb^�����U��k�O�C��Xjp�u��;�3_n�X>�k�3��s��<��+�5OӐS��g�^�-��N��(t�D��Ff/$b���X���0�8��*�/@{��)�79������3���Z�,Ǿ�kҵ��P?��5��JbG��xk>:�\�����.�v<w2%����Q(����Y|����5�B�A�F�{�����-+Xvh��лn��h(s�ZL5 |�]z����a�Y>�.�>�s���3}������U�x�@:������)��H�=A��V��U����h�F�5&�կ��{=�<L�����_ݎ��!�`h���~�7v
Ǽ�L�iS�"�~g�,���sC[���Àz��>�2�k3k��7%r����O]��i��� ��4R��.��n�]|X�bk�JY<{����R�^ЙO��E��"ɻ��V���Y��emB�,�ltkKDȬ~t�+���f�)�n
f�W�M�	8���q��V#	����F�7)���ӝJ��&	�א�:��E7	iOm&�A���8(����4_�[��J��Մ&�����N��� �1��+e2{~0���8'[ϴ2��4˲$˹yz㯍R�"`��+���ɘC��a|��"Y,���-���@@����===c���\݉LςI2��b�Omg�g7ݝG��3��8�;�`e�)���,y�_u7imZ�L+?��ۄ ����by�&�{��rM��Z���S��(CB��2L�AZ������oK�"@{K�:�ҾQ�:@;���8���{^��BZ ���-����oJ�ߺ"�	ӊm��
��k�iC�����3�k�B�`]�ˊ������Xޝ���U��9��?m����c�h$w�*�7MYF�5ϰ�΀�2Wn:H� �T�������2Gz?�ߣ~�j�Č����G�y��@��%���Tӝ?@%�4�� �Cr�c���#��	����nl=K��uwou��6�fB���=��*t��gy������I�	��N}�L�k��'M`!�,*7p�����^�N��O��K=f��c��)��M껆������6�^��=2>�㞺���+U�u*ew�z�$j|Եrܿ)G�qF���mf��ҍ�]�q[��8��	��u�t`��8Vyulx� �?�x��M�Ϩ>�N���9��5�O�Uؒ}��#6��)m?����ya��][�a1�u���Ӷ��cx�_�M�b]����^7���?�H7���9q�����{��o�#+���i���Qu҅���F�\�7��� ���z�1y�s~�js�4�*G�������������1�����"ϗ-��
|&�B��i���;�J蟩����~ '  �� ����������p�@~�1�d�ȩlr���@��b2wϠ���vGe�$�a��Û[�#�.��(���BiYI�x�Z�ި�nz���#� 
��IIK˭�*��n�kլ�LO���s'���(�	�ER�?_��9SUp���<�09VɍyY�\�NQ3E���;s�=<�J��6�,5������upt�Z1K�#��HϠ��z�l��j1����:�,�o �2�?:������df>�i5�;M�M��"Oګ5��͌��`�a ��*I�qP$$JTȲ�Z�[�B�B�7�xcw'�OalL�! �s��`,���z�@�:��G��C
PC��Kgt�X�A2�j�|���k�=��Ӭs�A�pU�P�
~���<��:t"3�y ?<P�[�U�W<��C�����M�u����bV�K�T,�b\+��!렝�N8�����6u��p�� ���&���De�&��_Y`�$#%)}� 
p���V��9�����8T��M�rY���g�v���W��Q�r��(�����1�Z�
�.�$bZ{�������O�٘J�=I)C��ǁ=A�� r�p����"��#}��p)�2�|=D5��i���|%��.I��j�<i؝���x��P0H����\�>�e��X�I��WI*�F�H�=�OL��*
L3'l�2����(���.��h|#-_t������/�{��u�"�5�]���`������=���������ߓs�~R�Lp:�^����8ȝ��f
��&6$�������P(}�(<�a:ԋ���<�-�^�z0X����C��)(d���^<�������_x1y	���z�tOy��w�_ݏ@�Hu<��)�������y���		<�n�����{ mۺ�^���;ϛ$��٘zu�)����d�zndD��m�+1!�؁�W	.�Hzi����S�i��R,���^��P1�pzZJR	����\��b]x�D���HL$@!�	�+����R�7!}�X�o�s���������H���j�~�[�m�j0�8:��L���㥟����{W�=�w�%���8;|��+��DE��Q���c_}�ΔQ�>��ߨ������^X��cx���MXV܇����f��Ⱥ|�b����Mh���X6���r�5}�/�!��a3,>a\��)=���e����3A6׽�6�ӣH�c��Wfɸ{��m0�\��������7�]a+-�l���*˻7����oll������
b^��^#��\e������X���cqy��J]�*s��[����0=�+�H�R�?F�7j�z�ZTr�(�>bh����3Z����4||a9����j/��b�&�xtO�H��=�'����!�[/1��z!?�,~�,xR��*ߊ�GF��X�'��4甍^m��J���tQ��x�t���L�pژK�=jw;N$��i�{se6�?�g�calޞ��l}�'ss��\�OEEƨ)�]�`�Hk���t�Z�6�$��9�uwSS�w3q� J�]�SǨ#�?e(F��r������z��'%�+|3�l^�2�k3����2ϡ�F�yG��Y�C�0_����*,] �b��aE����������~)G�-p�: ��A���[LP��1��ݯ�"7A�3U��б۞+�::Rx��Q�/��n}D1�j���,bݴ8���.��Zd��G�}c�&c9{�ρ���a�����԰�������vK�������6&�h\Xz�n #��*���\�I�t!-	BA���M����_/eu)N�"�����4�Q����}tv<�مX�0!�g�����<K�y=�I٣����jy0�q!
Jw���')(8��)�3q�PQ�N_V�C.h�yӛ���HK�����P�	}?����W���'�1T%��d��2
JJ�5gq���;��x�P�_re�VdnV�k�H�9�n��mO���gw�F!2q�^<.+K_,Nհ���c�>I��M<� �;6���������m�V��;`�Q��N+�d�0���5%����U�`�j���ۗHK����n��J�F@)�L��U=\��z��،���y�*����	P�t�ղ)�$%�`܂��;�$!��!`[KM�����kx8�R8�7JI*¸I�C�N�ZT�3���m&I��,���e��?4�7����@%�Tk/��N����!w�j�O��	"�-*"��/ �ډwV_�!b�}ɑ��#���gPG�j|e��|<sh�V_x4P�´���e�JR���m����!.���_���}$0�,e��kU��{U��ϊP3�^��\T���im��e(���M�!�\ʦ _t�Sd5'���N��T�� �E�K��jj�����S�|KT�n�E�'�D�rQ�y
�ڳb�7Y��Mu��
/�X�NI�(�`f���B]�	-[��D��zY'�Xm_`,	�̏v��;�����r�3���B�;�eS�q�:�D�~�\�([FX�>ԉQ�U����b(�G�G\���2�J��!�Bu80�U�*®IU��Qey���hA{���ʾ�ד��3��{�K<j��*ܭXm�%�U����1be�o�����z
hFă� Cޯ��3����JR�b��.vD��ϺPpk�J!����vn����1K��L7�bk�gY�	�P��Õ�2b���D�-��g�G�a���_��`��\��>b��x��b�5��H�B����Jz�zg2� XW��9�A�R�$�����x�v�8,�#g(�Ee-.I�_�D4^Y��
�9�� �����w���b�h�H��7R:�z_��jU��适Xo걪�E� ��pP�`�&5,ÖA��5�`k��9#YA�ɋG��*�9s�Z6񷇈�glo8��� ��؃Xm�;�6�z<?�Q-����g{_��2�
aԲ���ϲ��BRD�T�^��;�����K��Bf����K��Ǐ�0�R�kw�^�h�(S����1) ��{9�
�ڿZ��������ǭ��z�@�V��{��x���J��\�g��׊�t�d�.�<O���]�/O&j����z�t�0����Z6���n�ƿ�)� ���1$D˓�0�IA��C��^�N���7��i˪���R̵ͪ)דUW���s����(G�0��KO�����v;i�X��H�T��k�ZyD.�ynS���76ُ�j�~tٺS�@����p�;rb
~h&j�A���-̋�9���7�������w{�j���ƿ�j�_А�6y�$��\��d'��&|������1��4�«{�p�7���3�nJ6�^�l���\�v�忺^�W㿢q�qg~hh0:7^[c��i+�sM�(��7[������:p����"��(^v�c���⚿P��g>�`�{�?9��}������W�~��b�mapI��x���4��X��,Ql>��I�P��Pn�, �PӽƷ�����:Ѝ}�w|���L�5w�Hc8Ț8h^�Ie�x�.���SV�A�*�7冼��m� ��qy��n�KU���3���H��WTR!	9���ڵ�Q�F�ߡdP�S��<_����<��iS�[�8/{n��n�:5�\�R~"f��/z�~d��-�k�k��O�K:��L�r�k���5i�j���5eOeoN����h?e��S��1V���0�R�:�Ƕ[��y�|ڥm˺�I�yM��]i:�Բ��N�b#�����n�i@p�)qP�����TjP\�nU�F	I31���lU��)�hm��{����}�/VHώ��*�q����՘����x5��_7������'��;a�Q��1~XL���^u2� �8}�IS�M��;X�ժ�|!?�O�N[y�_ܘ)�A�������F&�9�i�1�ǂ��Xsێw�fs��^���E��k��ч�����
��ծJ,M��<��j���F��w��{���~2zo(���6}�=~�Ԟ�.b�y��,�,U�H�����9$�'�1Y�����%Ӱ�<�����0_	�$y���	?�(�_�MJ���㮒��%듟Z���3�"Ӓ���1@>e�%��_���.5ӎ�e��T�� �c�a��G=�
W�}��r�Q��Z�߹���+G����pq�B_W�e�2I�B���?U�jii��8�AA���:�P�Ǧ�iX:M�Bb�p<�G�>`�<s�0#���Q
��`�Z��MD+m$���"���'�?_�P��{FY>��ۤ]+�����t"�R�\S�z����7���A��� (Gb�uS݇�ľ/��T���v0`�ՙ�l��C�W�9c4�� ����{W&��+ɭ��Ȳ����yw$�i�~�W���N�a�����c�gE ��zX$~�36!X
uĽ3fN�3r׋z�����w��oi��T�\>��`b��)�77�70ԅ	~�1��Ζ�y��]�6��b��|���w�0M,��Z�������弼�O~7��q�p&��xkOq�d����c�T��:�b���_l���s7��I�c�V��VY��� @X��O0��?Ly�L�����]W�=���Ӷ�'V�A��#�o�8DEk����*��=+}An��_@�ϲ���~0����%����^5C��jGɠ?�6!����i��
C�.4.̸,wđ*Z�X';�J�O��f|�8�ryc��>���@��iRx�\m�Zz$��s���5l�0�wunk���{�3�����x�z��.�,A)��T�>���Q�I�)��?��b��㔐���0�m�~��t�F�Հ���@W^����(�w�x�qV�����D�\A)"�nF"#P	;��bρ=FM�;�=�^�?�p� ˧Q�G���dh�JQ���d2s6-z���q#9��}�r�i��ǽ�No/�=W�7TZ��ulԲ�%t�2:' $TEP���Řx'+�����d��sό/�ӱO��&<�@�I\�S��2f6�^��	����X��X�i��P�z��]i����4��&��E�PU|Ҷ�;Y��	w�=,�l�G�	��z�-�\��7H������g��!�[+�fU�I�z�i��w���T�ů����5{�2�7Y��jI�v2f8�1V�B���AJ�f����7�AM��ʀJ����{R�@������'@�l�,�L�=�p����B�Ѱ8��LV�x�k�$�U�W�g�b�[�$�өn��j��[�9�if��됬�﷘�ÖT��R��1��u|��1Vsa\S���.WvY���ͱ��k�nϿdk�Q�;_G��&VUa�۩4>w�Q�=��ߜ�S>W���m$Iz�	��3+�x�W�"���hD��fPc'O�� �)��[�Ap��DȡU�3��$�q�5J���Ck�_V�E���'m0d�nKi-͟<e��L�M�<����l1pL=��f�K���>�Lߚ߸|B�4��d��<F��.���=���ݻ��ˡv<��)��w&>o���_h4�bk[:��� ����O���T�:v�0��rJ!�'���J7�}ɰ#W��(�"�FY��eM�ִa`�}	p�������|�i�j���Z����X�xi�bA&Q��|��@�0�de5����C�4x�4t�o���\�-*�Q���@~�)��'<ܽ橝)���"��H�� 8��'G����ko� c�2�]��� K�7*�{�__�rW ]���XȣN��
�`�f��bW�;���m��	r���ܫ�VE��^-��>��j���n��3j��X����/�ݐV���2덫���)�y�ְ�Vr��2���|��V  ���D��EJ�U�M���ʈ�Ʌ�ڣtO>�7.~� 
ݐAo�}f��C�ܙ��&+ro������v���y���ck˩�sRW���c���s���&��$Aˤ,����W�ݏ��_c��/	^q9XX�ɯ=8�j&�l�D����]���/]�lע�#h`��XE�Ŀ<��c���t��pܝ���6U �'g�I9_`a��QVap�n��jJ�m�7{&�oo $���B�#O�E��d�Z6��;����J�[���6W(�b{ű����x�A�1>����� :�u2ǛLջ����y�N�S�wֈ8��ڃ@U�����Q���#��6g�r>E�u	ɿ��]��l�_�~����0F���/�zy������Zũ��{cB�	��K)�F�5��H��Xy#�h�\;xV�"�0��V\�O�A�z�J�":|��Ui�Iq�w	�г$�b� ��m�8'�G�?Y�?"�\��͈��yKj��,ZM���go��=%c�K��5�]��''���(ѥ�j$k�4������lːQϩ�673>@;R"��h��r��̠[?LU���ԋ�~e�q�^��˱����K�8��u���6�uj�f4�����г`�L�!�G�'�j�'����t�e�:��.!zb�*�F�|�r���?�}�A-�Y7��rK��QA����8�r�J~J�b昀��F���Zq�C�g�J �UhR�iMt�[7$��`-~�Aٔo��&�z��t����jjt�Q�iUA����&�)�t���S>C�����'��E��M+'s���"�!F�H��ۇs��<d��v.ҩ�+�(J&��LS5dG9_�;誠��J�-���v�W��Xo梨�;����x��Ix��w-���'{��	�m��p_{`,�Vlv��Z�/��J�&���+�� �7(���s��"�{���7	�{���x�{0EΏ#���E��y�l��4f����]��I�׃�қ�j�C��$�Ȝ�	����j��7� �J�ȡ����� ��Ƿ�9�"$�c5��9�X�y� �d	��d}B (o'ŚQ0��@u,$�ި
��~�Ҩ����^��Q}2j?yh �/����W�?^f�Q<��1��i`>�&� M3Nt �m�w1���
�	Ln�@0(l}n%�${�旤��*�X��W�:B̵L�h�l��r��6"m�︒ !���.뾺�}^6�'yB$��i���AoC����T3{;���j�4`�S�/���ʙִB��[JZ�L� �H�L��%�vѻ����~t o5"�^��!�!��n'�#�K�|췲bB����XjD������7az�+U�M=�?��] �L7�"���]}��,%ח �Ggs�P�������o?�ٟu(� ԛ_>NXO���S?��)����8b�N�뫤xG���o;i$�w��G<r�]����29L��<���P����z�9���Xi��C�ؚh�~�(ݱɢ��O`?5@�Y��n=d�Ϲ����:�x�|?��x��~��«�[^�9��F5(p6�^�dn"�����=�Ӛא�v�]�g��S��<�7'��ڝNW5D?,�ǋ�k9��Pn}aS.r�t�x7�vd�z��М�p��8�Aրl�C:p�c>���$~E�,u�l�i�3��Lf���~'�"��h�d5�Y��Ck`���A�I�ր��4���� '�����G�ݱ��C&��x �&�6I߫=�m�8�/0�l3ow�;��	�5S�5��5篽u��!�p�~ 8H��s��*F�V@�{�7Kq� Q�G����WIQ	��V��>5������n� ����������K���PR�Sf�.�'��E�T	���P�*:U��� �nAPr>RC���g_`r⭤����f]bL�E�B��t�\����<[C�N�F�����nI%(_Jf���-'Q��Hv+t���U��c9N�(�Ѭ<F��!��D�)�,z�$qQ�}��(l�H�����cr� �RS�V*Wx�� PK   ��dX� ���� 
� /   images/38cb4f51-bc72-4d24-b782-e5d855ce8001.png�|gX[n�c��"D���  M����t)���!�H�.���*��@@�tB(�	�����{�ϛ�<<g�^�]k�k���*�2�etMQAV�R	���"�˅�_������>��B Ǘ�*@@ �o�/Q���&�#���sGM�׎�/�MA���|�6�&/ߚ��ڛŭIЁ@�@���\�W&\]L��{Tw��_����(���i�m���?t]l���c���c}y0�"r��n>�~�2�4�܇���y���:]=�*���u:�����,V�;S8ܘ��`��������Q�x�_���YL�F���N�I���[̪��9���?-�%O�I��;�rv(Y�J�ӣ��7ǉN9.]^;sn���g��/~���7��w�矤��2�Oߒ�~f�s���&�`O�V��2������[�
�β�G�~�z,�x�T\�Bgv=�@�(��5������ЅM�9���<�T)V��m���q�X�
k����8k~Y�֖���Q=�AٗmYo� "�~A!�����K���WS���>�7��eO�r�D�ơW!ԁ����F�{�v�ٺI��G��h0ՙ]8jY����o�/8�\����q*���⩛6�萕t��嶋�Q��E����Ma��?|)�?�晬BuGQ¡S�wf0�'����򇞨�����?�����}oy�{x*��h����,���B�4�*���caH���%u<�@�a��%���{��PZ|g�$Ӑv��+�>F
Z|�[\�U��5���:��Gac���|�{I�5�݁(������Y"��S�ʨ)^Q/��β��抖��h��/�Jq�U�_��:\�K��I��\�pk�*	(���t��Rj_k��i�z8-o6"���<7��f$Rv?��&hD�K�ean��AO������5[�U�tB��&�lb5�53$f��K_�S�j�nl�C[A ���>��fQ��b9���	Ysl��^�䟧E	���"]`i�ePybГ�O��ݛqo���XZ�GXP��؂�J_�]�Mq&(O���������O��oW��4����L���T$mW̄��-�-��w�
S���<��f��p��)k���N�j)����s��y&D Z��!��5�G�D#=�g��B�*�kb�^m{b�R����P�xs�s=����� ���R^�j��)���h+�ݰ����oF��3q���#��W�Ev?��b#�Ќ�C^�,�U�4����2��A<�z!�P"Aѓ]���~#)Pz�:q���Z�z����A��Un���@W4������AK�WI��=�5���r@�+J�:e/_��&iК@om��*�2h��w�0*��;7(�#"p��{�갥LƇ����	ý�b����W���ވ��DA�?)^�k�d�\X0��;0�FM2�%/�u���go���ܖ�Yo�� BH B$�2E��o;���v�_9z�To��yK�b�mFrv����f��J ̴(CN�w-�)�zܞ�1�i�Z�3�i����Jl�Y�@,�Q�=�kI9�N:[�9Y�CznE=��ܓk�k]��l�q]G<�����T�D�P��@�[�I�қ̺��e|�������k����dr��r@�B��S�VIr%Պ:���B`�(�i���W�t@x�Dp�o�) ��jN���j���#��A�qN�U�8�cE�n68�S���3b�A�
;yTr�}�Ȏp�W�H,�j�b�#g3��)��`F/��qYh��i�/sD�/��kF)�h�4gy]h8�����q�Y��Mh&�$/)�j�7K�zpb�;˥�6��Q;���S�1�G<�?���ϣ I�I�4��t7����bn��:�q����6nDrvn�8�LVW=�0i�i�~��|�n'W�x<*�L�-2	6�eDZ�k���
c�@2�sŧ���#	.�X��c�X�;J����t�df�� �OS�U+��'�f��N�atn�ɒ�o"���
��Ū�A���"q�O�7z���5�:V}�>̐0�RB�@�
g����ӊ`2�9����L�fk@�R�wђ��B�z�_�04n";،K�N~�g��M-����?�?��8�Zo��U�~o��*yȩ�ʪ�#!���$���|I0f�g��
��[��W��s��t��a�rє��p��ӂ���a���z��ꅖ=��'`%�������^��2�	Z�)XKS��DS��U���LF��A��S�å�X�W�3����H���_�\�+x6�xN�3n&؃Z����Nշ08O|g�����L֪J����/~[0Th�r��T[���1�1�)?򥨧�D�RA��S�o
_�!Lv,���zk�21 ���~J_"�&�f�=S���Sw'�^�}�����lbm�ec	��=/�גU��T&�BK���+�t7���l��W��͡���D���,c
&]�=-����xUV̒� ��K�ˑ&0Wn��Ǖ��s ���*��� �f�I�$/�+p�{�T%�U��O]�&�d���i�\�yꉭ�9�-��"Zg	�*��dU-���Eh��oe'v�N
_��}d��g]0��c.~�R���H4_?�1sD����\EA'䢬�d�X=9�� g|�|��FDt�Q���6�B.ҥ:�w����ZZETyVͬ8��;:�s	0��hЋ����x��Q����8IR��<�Vv{t��Y?$�f���<�/
7���V���!D ��S�~�J�g[^����e/77 ����~�9��-�p��%!D	ܥ� �	FaYAwo��-��J1D6�	v�C�Ӓ�~�GP�(�m����W��m�rsr�S7#�MF��������yyy�ɋ�FjM��FK9˭�M��w'-SL�7B��_�/�.�<#��eRHG�8�(;� *h�B|��5g?���(�3�ȇ�'�;�8�>k0K
�L��1zI0���،��D�S�,O=F�;����T��-�9Z��n�]St�#�AB2��'��)ν����(S%��T���3M��k�U݋�5b�~VT�����4��e<4*%�\�㟣&,t��ds�ψ�]-�V0�r�����o�� �����SIb��Z�w��d������e�oie��bA���G̴�7>�=m_1�Y�yN�x����C٫��߿B����&�gP�<x4�
��OIIi��4�Xwk��u �<�W�_����C�-s��L�����xݣ�J>ս;��Vxhhcס7��v�N��������Q��L�ɿ"��٠$3'gGp��V��F�&Nl�-i��2,x�|w?i�6��v&D��S�O!hm���$�/|N=ӗف�ޤ$3�88 !\R'�j̀�K �L�">Q+�ZZN����1c3t��\}�������oIf�ۚeeeFIǎ�^;C�����!Bx���|Uz��P!�������%�*�ԙl����_���b�Ť?������1K1��f�f"����]�8�{�$��YW�K�aM$����C:�i�%!Ġ����n����ү]hi�Bլ�uBe)����w�rg��A����k��nP���ve�4w�.0WCU:cZ8����S�������inW�7���u����R�ʢRPd"'�;������ѯn��,�~�`Lf*����Ò7���
�n�l\`�GG���x��7=T��'�W�睘�S�q�B�ʥ�4�_^�5�E7����Y���0}�;r�C/v?�cY�5ag\��a��R(-T�4�������I���[k~�ͮ�<����a��I��Qx�����W!Vf>�{�mk����VlX���f��iz�K��x�x�ʣ;*��x2�t�����OK�� �뮥���N~d6	S<P>>;�3��!i��gj�5`�L�8��p���/:$!y�Fx��U�
�V�T�ZUB��F�w]�^�9��D� �OAqf�`����kג�����XN���f�Su��wW������N�� �#���z�wR�s�f���KC�ڿ��M3���z*���e�I"B�	"B�f�,�Sb�,�jsxHa���rJ����ؼ�^Kq�8\��>0�0��
�:̦x��`|q-! $·!��̨DO���_�R	�{	9��eſq6��b��܀��w�q����Ԗ��{��r(���a� C���M�Bk��y��Q��T�Z[�l�0�*�l;M��ٕii~^(�HY��<����n�0 n��U���@M�6!��$�_{�#2�8Z󃺑2K����6�R-�S #�h��s׹��cNqJa�q��]�q��@�2�� 3�.�\!ݽW
����T��^l�����8::�2�]\����u*��L&>�;u�{��zX`�����P������Ͷ��x�;ف|�V$�@}�ڲMq,3ǥ�ӓ���<�t�f�TދU��{�Lu�6Z��Fl�щ�&y[��V�_]=?�+�
��v����p�i��{�+�M-�h�.j�{���}�9���bO���z`D*��
�6>p���҄���3����+k@M;Z̔+��E�4��J,6NP|J������H�_dѤM:���Í!�����w�QO�z�>[��OK���i-	鳜��m�!�!���Z0�L>�O���V�	neD����[��.��zM:��H��9���9��Ri1�a��"�Q�
�s��<.���"���CX'�觟��	e���#gjٞ�+)���S�b+�!������<�ċ�b��^���񇾢M�E& �]����5�4i-P���

�W;-�4�R����㴂�S��l=�+dvÚ���\s6��!����L% 4��[z&�����tL����3�9�x�n��Ά?*�ڣ{Ժ��m�d:���Sл<+|q�v�N���r�� �w99������5`@0��	���uf��[��޾'o�g-����J���tk�Gp�� -���w��㞊za�_ T B�YQU���1�������#b!�y�PT/�F�u�X�q)�O�:ء�٫���3��}���`�;Ƞ�=&�pyt�\�0T��:Sx�d5-�BTƫ����t$��C�W;H|�wX���qWXZ�9YwC#�%-��]�6�]j%�3_�a�tN�[�k����j��Uo������,��!`=I%і������j�%���72~P���!��s������䚏��6���gW?y�u��7�δ��·{��Sg�̺�׸�%���P��!6����:�$���I��e��#@��p�N-�Ly�$Bd���5e����bY�#�>m<G'CR�m#�g��c���������㽺}�G'�w�dkm���Kܤ�U$AK�n8���"w�[+�;y�3=k��(�W-0���� �#���oe{�$�z<38?��Lm���-	��NS����U��%?=;����D�Ϲ\,3�
�-@�Cf����
VŰ�`+�3-�g����Y�=Ʊt��2I&����1�)���v���[��
U�f�g����R��UK�vӝ�@B�߉���n�u���ȷF�O����$�e2u��i�E���|lu�̥��l��.B�q�
d��	�Hň�x��f�Q�6L/@��T�?�]�K d'�����M����7�Ĭ����g��Y�/��7҇�����N����Ú�S&��*6�!c�=�Sx���k��n3g>_AZK1��l�eee��R�Dg~��U`�Xw��P(Ɂ�˪ȍ����������ְZ�����
5�ڵƜ�Yjj�$	k���7��{\'����6�Lu�T����E�4�K&��r-{��B;�u9�{b���D�b�C�)!���sYw��Rpp�)Xጕh4u~�P��i��L����';Xv������.'vv��3j)��&�\�dL�����J�o�f�t���ʌe�p�f\+C�+R.^�(�B%�U9���KĨKgf�d0?�;�d%iD5g����x��vs>����|n�����L��ӕk���̀����!C��G>�
g�#O�o���y����H��ȺEp�{PA.�Q�`3�-��������[v5H�������9Q�Z.>��z~����J_�%A�!?�>ڨ��y|w������$6"�1C�r$c�|+��z0b-g�Mo_��ᴗ�o
��v��[�C���Y�[����u�'�HxWٿ*S{�e�){������L�Z+X� ��}��UF�s���J��[(�Q8"mӪ�x�x���D�K��*��������&d+o׮ɯ0�8�R�J�따��c!�4�8}?Ai�m�R�@���|y4'%��ج�'-�����7��ܙ��T���l���r�/�Sr��6K�h���-P�L����׏�x+�e�׺h�n����ߟ��_�ش��h���Ӫ�d66S��|�h���UWu;v�`�JEN6�zen?�>2�gP;��GI���j���X*1�\�w)�^���zJ�<m�;*�>�΃��!��j���St�L{x�LZ��i!�Al����x��	�r"��I9�D��^�V��O�r�)��5��e�c'���W�p,�WUcF�=� c@�	m9�`*�'��4����=���y��;�c8�[�;	p@ۇf�=���@�'���jԼ\�8�l����椯�F4�Xi��H[��2D���ɶ!m��W���2P�B�Ѷ�17v�����6orԵo®L,O�l|lTS��W���R^�~튁��bB�~�3U[$Q^���+Dw�!���P�)�nr�}�bJ��[y"wʵ_˫ ��&��uJ�i��h6񻑤�I2#=]���f����X�z[���h	i�s}�.������9��]΍���_���4^f�)���]��ݲ�azx�%����#��Tb�;x�ǜ�.�՞��<lc=�?9�9�$�Ͻ 5Gn;���ɭd�>aN+�Xf̼����x�"M�Vq3i�GRN�h�rg0��2Xs3N�-��A[H�M�e�Z�S��/Euh���H r��Q�ﱌ�ҺG���]���SXe>řU�;����9J���L ���Bg�+��c�9KwGtӍ�>��?�e2�2�"�@��L��]2F���3�|aO�r��$���T�N�C|�/Q�K�����E+�0�C[9�W�*1K/����匿A�B8�~v=���K��B=�r�����*l�"�K�3Y1�^A,��?�y�9��p������.ƅ�ac�-�|DmN}�8]�X:������q{�)x�v����v�ID��jh����!uO "ge�_�X!+�V)��a���㏺
��%��&��/��m���i�j�|�<�cFl^��cr4�vJ`��8�Kz�`�B1��׮54�[�� `��E���?�'������=��F)ͤhf8A*\u�jq�WR�˜;pȂI���Ս�BA�x<�N1�P!I�km��*M�6��D�8)e��U����K̂������~�vV�����:�4�\-���_��J�v�Y.�Spk���Yh��:~ퟠ��9���%x]�\o~W�	̊gW^��b���x���`T9���R~�q�W��)���Xx/���u7Gu�RP1��ؑ� �`�aG�������=Е5�Ѥ�	�'�=���v����d��߮Z�x��\�G��f�L�����֫ޯR�&�ʫ�M�`a�� �@��/���^��f��iv풽N�c�0G�U\�h�&����S%�G�`�M@���j�-oa�-�I$'7���ml�� 4��ɋD�w�`�׎�O������n�C
��~�,�WE�[;j~�d�۟\�r�ؚ�O(5�!���)��|dɇyti�V� �$f�p��
� Ɖ�WF�2V�L�����9֖tw����u�=���JK_� %��F�'�WF'�i�ǂ�/�$G"�N��ڝC9hAe���=A�/znQj{鷯T��$P}���Q��]���v�Gȫ��������0~�����.?�F&�v��
������ÞE�aM⋌}��@�җc��sW�h$h2Vn���g��ɇe�p@:_@�IV�]ܚ֩�<�TX���Zg�l��xU�7�-�����:��H�m��u�U��^	o�����^�D�dT��<Lt��_�8����͆�mKb/da~�@WA��[S7�N����J�x���#h����=��i?�~�@��m�]᫝��ߕ�<�,�����o��t_�k����$@��f�в2�0G��~���^�xnH�k�`���K��vO��rk&P��2��s��[�	+)u���c�"2Y�����.c�Õ��٩u���2�*(gj-��������O���cf��T��wN9i1���ŵ�Q���eH�^u��P�\>�z��!�><���R<$��M�vu�0R��Nt+Tp�v!���)��+2$m^;4J{�c�j3�C���j��Ĥ%p�)�;*��*n&����pOԮ6��lA�������=����ncG�E�٢G\�9[!!Æ��G/���N��<~,W��E�fșjqp��D1�u�������g���*˺ć�-��Mf����?	r���B��g�K�ea���1�Ty#�e�����_��o.�|�8��bg�(̅� �<���m�wvv�?:�ז����6��� �z2�51S���*7`�&�̼�BK���r�]��a�z��� Gm$*X�_S�zJ���6sҨ�f)F}��7/��-x��h^�+�:'����lA2��wb��ݞ�]|�M�9eß}&�u��w�G].�D��j|�4u/��y��_i�ߝ�;`ۃ�ڜ�II��zR�O�:��K^�UnT�:�������m�~�9\����$�ԕ��$"���p��Y(<[S뤓6���H�������w���yyIXwv�0X{��<2E���������jǉL	F7O%���*�Z�G��/�H��}�(���8�q�le��!�7ݣђ'�z�6 v�O�Hv�-\�����&���(�u= #�8�ࠗ�Čz�X��t{�$Q��E�[���`P_�^w}�h녕����s���҄CjF`�r���]�Mm�l�/,��9��B�iu�'�)v�7�\�+�����zqO|Su��u��B�`��L��ںك��Ml.;Nk��a�uϤe�=�~>��t5�Î�p�.�sqҥ>���<��h�����[ɂk=�R�:A9��FUņ�>$iE<��)�,_���IA^;�#��):���c��e`q�&�@j�.��'�&ar��Bi��[y�����s��+H���F��B�/�w����$t�K8g��L�����rW����۫��G���f�M�O^j����K�]o�S�_�o��ʭ����K�!�g<�E¶��Ⱦ�%�cr'��/ʯ*kE��G7���I�(#��2���l�|�Z�_VJ]�wt�V�W��T���;�LFH�<�U�(��i�z}۰�;��tir���fŽVQ}ݵ=��`QY,�g�M�W�̑Ά%�{��r@2@�r���&��6���)������؇����_Ժꍿ�b�n�b����9�H��W���W}�%��!�R7V��C���/@�������2y"�R��F�'��VŃ�t�3˟th�@����%���p�"#�b��o=��t��
K��fW��4ț��i��6Y6^#b�=p	;*:?�]�;C��]}�`mB���t�%ⳎS6l�F��%�Z*�5|�8��N�]��z�Y�o�\o������x�� ��b�U\�Z�w���3��K?���t����1d��E|�d4b�j�b�.���M2�1���8�<ha���^TU�/�
`�����#^�>ͣ8TX�*ג����K� �ێ,��/��$!Y�"I�!ʽB�Ъ���l%b�l%�Q����F)0%,����������- 13�7���|X1���^Ϯ����z���^I�=I�n�\��nU�2�~i����@@�VC�O~��&����@��0^d���w1�e�L=N-]��*?�0�ڪ7��艧c�"sT��'�a�wY�1a��^w����+��?(�G[��l%,�P��qmV���m�-��DWWך|���5�~/�՚���%9�Z���8҂��ۻĮ:K>�'Q�� ['(a�����������u��)�No���ɜ�
L�v]��ߔ���Z�K\?��@����q��U��۸�G�ѡ��.��;��rZc|��em��ж�1Q�R�O���u�؂�y�*W��Z��3�
aP�ڻbD�5����<:�_�G~;xϠ�e�ct�ϩ9�N��))��LA�mT�#��@�gW����xI�y�� ƂH9�U���}#�v6���שp��$���((�17ih8��B�E-����K_��,mVC	��
������k���.EA>�F�Kq1 wJ����\8�K3Bg��������p��|�'��j������ݣC�LGˤ��U����C�܀Yvd�����p�GO�L��y��,D%�UĊ3���쁼b����J�rL�--S��u<�t�=��m�{�v)^@�7��X�}0�z������hF"�Jkz϶��b*�N�]�X�������v���ݯ䇵j:]�b�0�L��h� �8���Id�����t��㒤6]��#���v,6������i�k�\�,}"h8��6a��d�k{�1��?t��������m���o������J��u�^YK����;���I��@2���I���>~��ΐ�*��^@�ˇ��
B Pd����Qypy*��Ip�j��6���7��t�r���Wx5�쑐}E���}@v���(XO���_�T�J[}_��Oz2h"HR@��.��>*ً� 7�Z��Z,	YK�$�2W`n���ɈJ�t�56���&I�B��]4�z����ᾭ�q�'vc��j����<7�T	+�=��^F(��s��i�p�pu��M ��w!�QC�%�{�(�ӏ5��Ǧ���%�-jĺ����~��>��J�;���=K�@^cč����I��g_�^���za	e�jwn��� �A�
�k�G�F]E�A�m��j�b��[e4��b��C�Οl���#���p(a�}g�$ ��6/���1�(mX�5��}����u�g��l�0�t��y��3Y�(o��|,`��������jqT�n�N��;�v�s�'�N#-���Q�m\͞�Im�]�ID��/�!P�{;��i�:�R3 ��������$Z-0�֯�X��Z���\�@��$z���u ;E�լ �m]M���F}bZ?LV�C=Ji�/�m�q���r�u���̈́���	*���0���
���4�?��j9�î�y�KU�2�uȗ��V,!�A��hxx[ʭ_ήqH�5�a
&q�ɇ���^������M'ܳ�}�T'�D�ԎI{&@������l/��G���a�WR�cPC���²N:�\�f�5��)e�n�\v[�ս�~�n_b}՛���W�Խ-��z-�}������`���3�"�J.m+4y惡����/`έ�@�D�
��X�B
��uԯ������)$ԅ��X�^w����#�<�I�Sꔾ��h� �B���)�.Qy"�F�Q���L�{t�ژ�G�]�I��`3stT�d�^�V�!�
�7��V��3��T�<<9
/��<LC�,��kr���'�Y��ܿ���ѕ��4B� ���,5΃@i��ūp-��bSh9�n���
�l�ԪNA�����2#9��e�M*����kX�n �2��`���nT䚽�c׸?��@&�QW�nǳ�Y��%]ʵV�=�4��ٕ\�k{�`M�o"o:x8�0y�eg�پ�2��Y��`�5/kMŒ&���B��p�?�sN!J"ꎐ��=Q���9O��]��s):�IB����\P܃67cU�E~gk��Ӛ+V�ϿdCK�+iTYl4���Aԅ�І�]:��}����+���㈆y		4��R���^�T����ǖ�d�Q-F����������3$�\��o�j-���.��\W�D%9�u�4x�n �ݰ��Rxtչ����E�� M�#L����R@d�B�r�k��5���J�2�OY�`M;#����#?!�o�x]�_��:2�@יv���ܓ�__E����v��[��E�O��2���z�܄��0\V��Mk�άap�9h�-_���c��m��F&�yl1K�XMIL���kuV� �rJ3���G�R8�YZ�m�< E�F��K}7�X|��af#�W�i��Z�Ɋ�/6� wsf���w�kP�W�Q�f��0�9��=���h�eH��Q~�%�����ǵ>�7�Ӽg-�<��BB�.G|:y{�޶���p\��P"�d��~Z�,�z��ե#E/V����s�v�M�5D��"o�N��a�;v��}����~3S�n���{�X
[�Æ}_eu����Vy���.����TH>�=��r.��t�ut��W~(bX	p���|S�u�FH/iL�/��a��-��?�E�eY��&���d֎��Y@��a�K�0��{�uF��Y�����R����2���H0]/�c���*6���	̴�������������n M�2�O3߄��Bl�2�n��k\��vp�-z�~_�>)*����)��I��[��'�߷軧x�?�y���g/���wMVA�v]2Èg*u��.����6F���3�W����+$j�mWrR�[	gpq	�F߹�O]�[м�"K~8�|�.�:c?M�]J�9-<��7�R�kZ���l����DK����s��1��佴�*��v�ϲ�8�1�ͅ�g� -���<����7�2f\�هQk�F�M֡F�U��F�S*
P�d��I�V��|�J��i返���@�ؐ+f��^#1&4%�;�ŝۛ��1@a1k�vV�G�b��݉�wGR�>F�F\h,���R,�>F 1����ja�����o����͜��0��D�&��0������6Y!j[�dP�#�sV[)��i���`�x�b�����P�Xr\�/��谖��G��3|5�_��{QONn�, �K�d�+�˶�M�)��L�7��b�S1?~��@�o	����m�ҷf] ���J�o����H|�19\x�ڜ��5_���*��IQSS[�~\���W��)��Q�������o���I��O�*��R\T����E٨\Z;	;��3q	��*��q��Xѩ��xB�x�>�sq�B��o��}��{N��+I<��#�+s ~wz;�>�����T1�~��bf������کj���ZC?���^���j�.������	��S0O���G��*��\]u]�U�MJ 36=���IK���Y��a�Sj�Ϙ@�L��	��Q��7�'���Θ�"���l�� D��(n����3RY�����l=S�%7�k���X���2L�@��X%�;"��"$l?��0d��
$V�۲��t���\�V���yTlo�%D����� ��D����m��R��!lg���lz�����}��U���>�	�9W��.����<��� P3�g������Z�a�*J�F���n�K���gq�m�aX�����T�����c���4W����j+_��I��#���x�6w彣�����W�c�m��ū��<ϰ㬨�t�\;��W����@�r*�
2������#Zؔ��[���Ԧ^B^��[�V����Wq����N}�I˛��d:)Ǭ������RD/-��6T;��p�ro�nsm$YE(@AD��ob���ͺ�`[��ؗ�& c/!0(4����f�&	,E 	)�{y�X���	3�OU}����`�V$vGtjk[�[�.�Q�s��B�MhL*��W�pr*���3�k���𯆀���;�\�y�����_f�Y�3l&@���_+d齎-H��3�2q�iA����q�]�9J�V��#�@�r�\��DjuݑV���WZ�[�b�$g��J�I���aO2��<��F�||�I#�T�Z;�x�����`�zP3Y/����1b��D��;��&�dC��9�W�<�V�󍾆ZH�w��ƨ��<I�~��,)��Ҍ�8%:[+5<�g�6�u��5_8��)::��Q� ����?D������C��m���]��s�^�^k2�@�-�i���$��x�g��CB�U@(��29�W��;�;o4q�V�m��$�y��i{�ٻ�����{s�YCm�'�5&�7�)�;6���L$6�ܑ�����d��UH��'�A�Z,���n��iF�ݖ'��|)��`�x�$*�u�?__��x�'�n��Wq`��$�(��Cxk�<�\�6�������w���O�Ņ�e�ЙyL&�>�3_��� t�.w�g(���z�-z ��>c)q�}��YL��ǏN�P����U���Ɏ�[5�5H�d����j���0F�Hw��xRb\��6`R����h�����m,���d�a���7�t�؎qCn���e��=�b˵ä 2�BU��[7�"p��g�'S��zo0}W���eI'�LS,�Zܻ����8������A��p�#�|.f�2���ñ�r��5�u9�3}�M���3�|���X��̵��n�Zv��g(ǔ�]͚K;��V{2.(��F���镵��%�0�nR���LǕ�a�H����=*�V�?9y�������?�a{r#*�:�!��'J���H�А����׌T@�y��
����ٛ�<�Y\'����-�F]�r�?i��~�?A0�/��멡�!���KW��t��d�K-�o�Ʊ���Ά��lSQ�k��n�E�I�J�BB���:|�^��=� �D��J%H�S�(�Y�*p�Hfq��`��z��{��n�Yl�MT</<|��I����5dt��ﰇu/^*B��Dnǚ��[T���p�,n�koP�
��[�Q8D�����p-�qV��vyO�}����v��E���o�
��S@a�;���[�3Ln]�p1�Y�Yt|��[�7
�����ɤXI`�w�Ĝ�#_���tb1 ����|�NU�Rp���9�qo�����O����E�D�+��!�?�ޒ|<Ϡ*�d�dm�#��!���-y�\�?ފ�F4�S���&e.������D|G�Ą�M ���S����Ы�����{d	��a
O�����	��F�Yy���@aA���k�9�m\F�KW���z�%#)����9�R�XF�^l��t�E�����Tm��d�|���@7qЭ���U2�A��u����2O.�mNտϔ9�v��U�q"֊(��Ξ��/�[� �"��ٴc�"�Ȼ��t��� 1�l�bs���/\9��kN��BH�%���.�J2�\��i�q!�4/*y���W`��]j����_��>{��pd����g�+���tC_�Em��X�W��&uAA�W���ɓwR,��R����L�R!�)cQV�| ���$�] ��T4xo粰j?�����݅3ʕ�Yǩz?����.�ru��$�=����]r�ѸGmPl�b�*�f
fN/�v*�#��m��Sx�\�p���3uL��$jkA%���ע�� ���;+�wA�V� �<�=hU!oX�EF�;�2|8���	J&�������yL�a4����wE8�N9�B�2G�@8�<�Ը���u���/�z7 � �4�Y�&��{i�b�B�|�XN�cÑ�	��^�	�g��F�tJ^�
�ѹٱ�Z����[�Q6��>2.�od�����,W�r�{�C�����t��:5OO.����_R�ޝ��x�޳<��D�S~�9��AJ㺷w#^	|�P�ՠ���<)�E�H���x�S^�2�v�b��lW/�V��rK������E�u's�d�_��eٵ\����4-����x��Q�	�һ�C�C�{�"����S�Ao�����<O�3�]o�-��w���7�r;.$2�O`W�A�-H���������-?���"�#��	W���8楙�̉{����OyQ�Rn\�����4o���5�j�b3zu����u�D�9���PEa�b�2�3C��Jjb�^7�|w�/�(S��de�$�{�^c=Pg�Q��c�ys��I� G`��\y�9����3�\g�%�^T��ܫ ��u!}� 0��37�=0���p2m�~+��n-1��KT��=�a'�FP\-�v�pZi1��pt����j����7�b���������"����x���j_��!h(]��3O�D�F�O��f������{7;(8�w���ȍ�����'� ����Fr�&�H�����#��k�=2��rb3�����|���G������]:f��0Z�)�-ve�2��*Y�ŐCѾt���b��f.�/rk��}lN�]�Ȱ�l�˻�2I�wi��z&c :x�H2eW^x�+���p���.���.�_K��������ۋ0��|��}��
��u���>�)1����/�QO��@w*�Aު����Fd~7BV�4�گ����*=�6�Ƹ"^x��ǻ2w{���{���r/���m�W�9��ӎ�[�G�Ӭ�Po5 �����Q^;,�<�;�7#j�$�#�Ck���L��r��[F� ��Q��.��z������j# ����� ��DRnw�k'N�F �'�UA��.>���.Øn��eo^�ɓi`Fm��?�o�Hw��&� ��~��y���:8�V|N
�d�ȯӲao����}�&e�Q���]!�5@�[@Ω��"��b%���}K��Y>��˿�`�[�2�9�2Yh�I�W�"�Dޓ_%�5(y�<�޿�"���k���H���j�0��e�V�[q�&�ʣ���k��T�JL����q���X���gUd6�uGj@�W�{�0穡-�������t�Ɲ���ُb�p�֤tDѼ�},�J��nT�6��Y˂�<=D����ً�4�"`��a>�ǔ�T䢀v��ϼ���6���FQC�o ��_�L�<����F,���O����) �y��y[ R���C�=��[���W8=�VE����W�5�vac *e!�� ����n&��c�0T�{���ݠ"  9z��c�t���=����}�|�����\��+@��}�	�،�� ������9�V��������/,��i
/-9�̚�������sMhL��QR?i�2"���<�e��>���;�/�VH��,E�U�c^�ΫA�.��W��O��ԩg�F[�{[�xVh�`Y�>
�]�����%��GXk�]�2�//�~{�S
	�{]$x�e�X�|��y���^��!����oa��˹�	�^�?e��5ݰ5x��|���ʹ#WS�\jU�p�i�"�=�"⺎v�`Q�N|0/u�ad�}j���/�l�~�HBm�bu��n��&� ����lo�� r�+�	��w�_\��IS�e�z>�A�֖ B_$P[ڠ ��@�6J��|uc����?�5X?���X!�$��˚I�l��AM���k�)3y_�#l��{[v׸;Ao3f��;;��ٶ��|�^IPs1�\͓�H��k\�Z�cU���[��!��4��lqB�_�� ��P������;��Ϸ�j���ګ6_���[�_�(g���A[�vKVl��Nz��g(�릋Lm���%����bD�I����g=YsL#�\�,�l=ȱ����J������6�9��ܣ,������sq�r &`� ��4+��\ӳ�F�q2��U��m\���B�۟?��r~�dKW�jBb�Qj��򃶻��tr�I�WT@@JL�|>ب?\#�{�X��6? n�F�$��f;��� ��������d�����=�{�#OWv4��D	"���γ��nG� à�6��o��3���=F�$3��\��[/��	_�U:��Ơ`���G��9K۔'a���#=�=xA���j�eJ��~� :���&��+�=�����'�W"��Y����Qx��Vٗ�<�o@�rO���@��$`����c��L������v,f�o�>���":�}y@��m�����癁m!4nD�je�4�O<�����PN����e��B5�z?!�d,TSdwHNV���pF�Q�{���t���u9��a;΃:���X��RR]S�\��A �?{u��2��{�������\e���wx)���:��5��HH�xC}U<W⻗#˶; ��[|,�����9ZȔH�r���������X;0����R���7��;��9�e$d��>��ޡ����o�c9���& XP?G��9�H��bqt���3=/�2�[N�3.G��Cl�w4O��8���"G�5^�]<[�#���9����֤`�a�/�����t���彔��°u���ް��(,����鬵���1�7�3�j��,��~δ�:��R˕r�(��J���\�ǈ��v3��/K��a����FN�w�χ��:�{-L������!f�srC�֪�ߕZ	Tگ��7�O���~�Ё
n�Л����� ����?KI���1S0l.Lt=@��Y�� �QF�?]��E㺦��n����t�v�nxn'�-�y������"�|���w^;�GGof�g�f��3�Ys�ٹvv���l���dL�d@��5�aIپb�_m�wg�`:i[�}� h���Yv�5����zx���Y ��l�Pf䦦���ݥ�Rx����{���s��sn�}��rc��yO���}�hs�S�E���%W�ўOv	�H��,�4����{{9�X�{)/G�g9����amQ�иe�{�Æ����Ꮃ�v�ߏU�D9�J�^�Hdl��B�8��ˀ@$k������b��5]a������O(���q�T	�i�vLIiI��T	s�T_;�
��~�|e;K~�!$��d���s�������s��.��y.���zAe�M7�=T՛�O��~�����
w�f���ɨ{^3R2�+��
+�	��I	"JZP����9��rg���2����mN��3JՋ/�n�g���5��GT�0}�п\&�"��8׈	�;�E8�f�Oq;��^���
A\��]pq���^c��σ	��/�̖���Om��2u>�oT�_���v� ���)]�p���nn>M['�� !��!+�l^��ъy#�~Y~��gw(j��8
��I����!f?$���\aÏ�*�ru
�vvV*щ��Q���0PPK��CʭO��P���K�w�Ú�� ��-�Z��G>j���	�)+�������Cju:�	��aA"�l7�^Z*"���V��w',c���b���_�:�������U��n���˻��N�k'h|/�G�\�F�"�2��!9��O����*"\;�'��eh��ؚ�GE�X���W��r��;�VW�UlUZbt�dEbQ9n����{��R>�_�
�#ٱ��'�	��؆_��gpG�ǯG��'G��:j��cj���4R���I��'c�J �K�>��Mٝ���j��y�I�e�7o�b%�K+r��.�n�4���9̘~����иE<�[��ą?��Bs>;�A���(�#��ݧ��!O�����-@g�d�Bn����4��H�;-]�{�������=��� Λ��E�F�8�aOާŰ����v��#�ꗃ��]Zc�:�k4�P�a�Ms����VC�����S*'+g������x�b_�l��������pFP�]/	:d�-x�F>g��!E������1A(/��Ѡ���#�L��A6�թ���ڼρ��wD�S�� Wԍ)Vf�Pܢ*��[��v�R3���������6u�#�V:�o?��P@�j��!��j�՟�5�7	�ڴL���<�!J.r&���|\�y�	�'g�vhu�R,��K��g�kN������J��J�d�Y�.��/��;z�w`t�b���R��`�P�E
�]l��9�Ӂq탮�,����*!�'�� �O������!�C�Y��(�m���q�����	��"f�_��L
d�Ch�����g{�oVV��"�0��z!����i��;5������&r�զy�OTy�d��b'zuc8�:�<Rc�F�A�A�j�4~����9*��[��VH�N#L��j(�MӽM��K�rm�Ӏ�Ms=��|��DF�)&�"��ϕi�6
6�E`
f��[��R/�D�մ2DI��ߪ�db�������;6�ލw���.vdaS:d�P+|	��YɃF��R�cO�4��9&)��4)��v����7�	?7�JR���>PNy�O1�[�^nog�ɷ��t%� $}n;��{��(\B�҈n��8`Y=1�۟㝡Wa�MO5_����]��2Z�w�������`��\�Ʊ�鐑�a�i�J��0���$��N~t��g>"��~�����T1a�h��}\�4�S�>�������3r�m��*�OA&_�iq>x!g���%Q/�u�ؔ�Cx��a%�����ira�2.YAS^�U�l�?���V[�'�~|����F�C�����,մ�U�W�7s��>���{Mi��5Z�:�=}��m�0���莙��ߊ�Y�e�6D���әq���ݩ]A1�e��i�e����&=��lmn�5�KU�3.��8O�2�' cU'����oU?l�G9��!��Y�D/Rs�ot�N�y��۟���^�6��L&ߨ�֋���YG���ˀ+�{��9ޅ����O���,�|D!����˥�^�~�Qn�)*��\�CY�8O�/\ԃ)K2 �����1_�R����g���7�����\��M�vZ�JJ��j߷��
������x�@�W�٢G�����*��{h5#%�fͫ���&!���;�0��{��T���F�Jځ��qp�ßc�&M[�k�Ӎ�0Cvy*�I&&�u�_�m�'�ήW����������buJ�}�D�Vݶ+9�A�En@��y�:]T��DXE̻�RFj:!Xt�4����z��|aGC�������
w*��t�N����$���ɜ��f̶��� �O�j�-����rSE��oc|`�9[� �?���v�*�Ѳ݁�6���Z"x%����߳ T����"_���|��9L��a_i�e�Z�&e�aXUq�8[�p�����M�z�-Q�䔪g�go���j`�Q4����������oh��t���w�Fv0�����3���tHu�)�$]��"�\�m{�Ź^_='F��R}(�A��et�J^��)��oW꿘4)�@��q6G�[��ʮ�&�	���o*;m�V،%�^�iB�o��y)�1@l]v |'8��gs�����{�;5e���ea�!$��Tb�t�b?aF��W3�V�]D$���R2f��x�Ú�ml���������>�T"2.�����Hc�$D����}��
�z���l�k�@%�����a�,3���D/�x�|=D���&nڋi�:6Ǧt�Ҋ?[-j����ۖb�'�2���	�]塳;��}�;��:'�k�L��!�[�
��$��>�?�_�=�ٌ�;����ML,>�����1�|�W^�KN�	��+��e�
�E/�̀$�3$�*�y��׋��9ާI�g߸:���������r=2�a�oe'm�g$�t]C/Ul�h��48/��T�>����d���$�(�y�yvQk~ş=��2A���v c��?��?�j�O �:Z�ތ�:	�s4�Fl��q�����G�>*��Ns���7�v\څƵ++h��J;�'��wΆil�_I�O{e�MĊ�Kr�6�����#���^L��g�&���,e_��b�%o&F{9�z��O��+�a̰�q�}�r	�������~��/)\˒���ɞ�Ϛya�n����񭰍m��}��)\����%�&����a��g�w|��\�)�L���;w���z��|Ϻ����n@�ȺՏ�fvzҳX����V�CI��=Z̠��)Si�$�W	C�ɿ�?`�ۘ��.s({ob ���c����E�����m���w0��@�;�@k�x$ָ"�Xa�i�R,ee<0>��%�l|�yw
B�s�Z�=|���W�Pۉ��Y��ɿ�3L����3ū��N������vP���'����6�kT���uYeM��O�K_�ޕVn@>�z�uMc�)V�38_�N��t�Y�.F�p1��
#kbފ���{�-����x���>vw�H� $���QU�T4��>�����x^-���?&／nЭ�� ��&6j����S���\�������d�<�F~������4��e�����9��ƐC�奴�]�AJ�|��nۑ*��}�_�S�K�X0oYV%�35���&lJ8\�J�݁�w}Ao��
L�� ]����u�fx�o�P☺�����j��44�@ڕ4٧ݩ"�3૦8F˧>��E�|��� \��V����+�*5\mٸ�o�fg�`R�}}���B*0���+�O��n�pN��e��rb@��u����KgT�} �o􎊀Y�E�l���es���I��)]6�P�PY6�SxS���L��Л�����o~�x1��O<@�{��ߥ���"}1LJhB����"z�#�c� 
�{�|�e��uh��e\�FA��O,�n�=�?��ܵ阬!_�mtn$��.�QDuX��B�j+�o�{O�Ǚh�V���(�V��b�b��K�p&�J�5g�
��(.Gϝ�,�]e�� \�v"N��[g\כq��G���2�
��+�U�o�b�����ة�a��S���Gϓ�ZA�K}B�A�lw��Lp{k" ��@ᭆ�I��f��C�
H���ˠ��'ֆ����IܶwIF�@V�����6<c��7:�������(�������:����Gg�Oܓ/��ɶ��cb�h|��x�>r����Փb��+e�P����#�d�i��=?�s�(�v��]������o������h����W�z�t��P�`Q_�����/�޼�#�wl��*���5N��f*�RA���c��\Yo�3U�q��U�(hY����յ]z���1�
���&�+��ԃ�#"}�i���Wl۾u�s���[t�{�5�8W���)7����J����΄kjǩ�%R����Zi���j�%*��f��y��?)�n��:)=�]�>e䤫��.�N���1V�=�x�t�i�2�)�S4�04x�hԾ��`?�XoNG-�Tݍ)�����V���ՊnC�#�V��ķܼEk
�0��q����xF�U&�H���N��u [f��zK_G�Z�ڮy�zEd0#U�Z֠�K�oe	�f��lr�����9��@�;�k���1qL{��FL���������g���#.�Y��2������g# p )�&U�ht�t�ns� ���wِ�+�٧�o�j��!)�l���G�F�>��o[�+RQQɔ�hj���hw�Ym@t������޺g�}���qZ��
N��7b��O�Z�������,�FXW:J6�AB'�{���j�@p��}�U7_�.�U���Y��^�p~��5����`�#�nm^�J�\�\�^K�B�zs(�����w��K���yJ��>=��ʅ����
:��m���N��:o��Iz�"B�b\.{,٪7ҽ��w�\�	���5����tQ�Ȫ̬�+M��0\�'�TE��[��M�-��~R����9�2V��$�\w�nq���q�v>�����y˪zz��K_�]�g��'S�̶�M�NJ�3��4� �ͪ�OR�Tͬ�����L�Y�W�a�e�M��֔W������Z$���
�
����O�/b�]��\����77�JL|�\q(y�Q���K���t�V�6�Ě,L�{���T�M��M;���.�	qsJ�"��O�9���^�|D���oט��<c�|��t܍�I��8>�h�U�U����uLl7��ѓ��3i��E�C@�qC��7y%TнmO�f|�}��K���lƮ�	��DDQS�&� 
����v�R�5�~���)�bu�������T���'?���9��~�#��į��/}f�@:�-did�[8�.!����]G����߱(����Ր�(�>�I������EO�h�lI+�fz�T��K�V�?}j�ZJ�� ��{E�b��ӈ]L�����ֱ݈3w��N�u���h���V�,	�H�b˼�-d�gHe%�l%�)ò׈���������E��L�cJW��U��K
s�tlygggtor�?��XNDAl����F'���_���|�A-c�c�;T�k�p��J057'0��מ^�����qF4�n����Z�gx��,�ƲQ�bSvH�r	/o2~-��t��%�>dӹ��i�����^�b1��*�v���VӔx�\���d Ӂ�������$�'lm}c��saIT9DL�	h�*�77�#q�����r��-GS�����N�z�n����3�����1�v�E�G�sU������(����w�5G���{o�����^{X�ܷ`�MOΩ���$ w�Nx��wI�egI�T白�+	�P���u��<ʋ�x�1���VV,b�r��wtX��0<��G������^_S�af)��Y�<�����E_`^��J��6@��v�k4��,�F^���n���� �?��mCEA�2�N45Vc]�%���N�Q�*&3K��?3��������>��1�(}���n*�6*�c!����t�\e��k���D��^2����=Y�t���"�oRVO�CB�p�����l�����*�V9���^Ot�̪Kq��7C[�OF�D)˳��*:�E���cRߘ�
+ɝ���>�hxN�Io�?�L�p��'�硂X��N ����T~o�s��&��ț���)M^kȰd�i��W������ޯ��W&�X�yi�sy)L�.a�Y�պ�;m|'p5��"*G��4�޴-"�K�q"�����a����W�X�SU)F���������(Ժ�u�@��6�/�$yZ��_J=|1M�qp��Ūz�����^-G]���8A���V(�� /Y���*��N�����ʲ�Z�_Q�1��"w������E-��ŲgW�A4a�ّ�se"���[cK!.��m��Uv�~�eֶӮ׈-ߣn<_�Ԋ�}�w�&�Z��ƘVޞǜ�l�n��l��.�H$���|Ԍ��6q_h����g��Ɲc:
+���\�aE�Sxfu�����w��i��Y����3dy��@ ��ly�n^��ai"#�6��}����N�d��!]2i:�ĭ*�ng��醇�:N�,igrfr,���u?oʹ�������=�85m��P����o,hZ^Ӵ@ӫ<��4����=�`���_�Ϧ������O��1Ѯ�꾘ir�����\��O����ߖu֨����i����_}�3تbFg�ɏ���/2ɨ�� �C7����xiz���o�3���[����Y�6����Uq��)�U /0;4��m�O/�..�L��b�6
>R
f�}1M����q�=FHsj��'Dt�͛A��`�3��������z���9���H�C���)�� (�6�B���m��ھ4R9~�M�ylO�h�6���4lh��ms)��Tm�z�I�$�}�G�0������A�Ұ�br�I�4�/�wvj�5Zxly��?�=n�E�Qj�8��~�g&%�8���SOI����,j�/��Դ�M�k��h���t6r	{��?T/�կ�/k(i�V|4�t���qx���4���a��X�/[�ko�
����C݊���!�����x8����A?�{�y��y�� ���^�G��d6T|�f��c�����pt��;���j�07'��C���٢i�Į�Wv��QC�٪	�c�W�͉i���I!�}e2�{+�EL���B<Z�j�e��]L�^�,��zw�:ܽk�cZ�%�핮-'������[�h�n�SuCnB�o�j>֑s����،�Rv[U�����>�V�b��-/,y�?Ø�z��f羥a^�rÙM;�/5��W�Ж�	<�>f-9a�~v.��&,�Es� W��1�������x< ��&�)F�P����i�*N"���p��<�\BB�n��p �ԮaM��w�cf��&���4���=>��?O�V�T)��A� ����;@�DN1�kF��Ʉ��$���� 6 /vH��G�V�;�����s�;g]Q����L��w]� kW	�Q�D4& ���`]�Ԗ��=��t;��έ�y_�~�ݺ��c���c_���hY0�K�"���H�Elʝu�c��z���#}b:+H�/C�?��a�r}W	��>U��݄�jS����|�"�~��|�?t�{��E�����q��u��t��|fUZ�Tσ��u~'����^ x��\�@2K�������+ ������n�8>�|�dP��:��f9ejX�

Sܭ�U(�j���͛�Q��G��M����&�#��.��]5���['��$,�_�a�I�F$�����۫�c�XWM���Y�j�1��"��K�.�^���@X�߽�C/27��kc9�l:��e�s��(��P3���{�}��٣���g?Q�
'U��1�m��\�{6�ҕ7�=P��:�N�51ǪX:O���Ku���%Y�츍\ ,�:r��5H�iJ`\_z;\ޫ�H(+����s&I
y�(����q��{��r���SS<�K��TS���?c]�ö�zWPLW��B�x�J���8�$vs�}=q\�1ӛ��g։��m�5�.r?d(���}���x�/^�ԕ,�.{��_���b`�q�����a�J��8A�����mk�`���7Uɋ�a �Ș��a��l9�=w~ϙI_�#�I6���뭬j�"5���z�5Z��ZWY�@�d �Ķ���7ih�%�"2H�#`����C@�9�=�nm��v�4�F'��̙[|��>vB�xM�f��&
�t�<1>�rHl���Ŝ�������m��FgKp�~�"Zm��{�l�-v�e�}��/%���n�H�s�I�~HuR=��ӷi>@g�^As�^*��	*ϟ���	b8��/�fVw<�e��=�b��z �����ķE@ߟ�**n�e�ZNLVҿX�ݷ� r{ ة���H%��씌0�^���E�����У�%׿�Wڰ�:-���l�����Y����h
�4r_N����ϛ[����ʋ#�;Х���<�F�.�ܜ�OM�]E��[���}y��TP����Ĳ�9�K�_	="R5ap���R��&���y�qi��Y��n/��F��у�s��G0��Dye�e�[��TMqd[���V���+��D<-@\��(��Id�&N��.�B��j��]ʚ����-cs=��Mn�i[?�o�Mȷ۱2a�\y������rJ�^���3���m��AQ["򗂧��?��A�T�T���{�S�0�Ŋժ�w�啠X�Wv�Q�wZ�r�Ne-�b0���!W�����?;}lmfc15��o����Lѯ6�"���`<��VT]��L}M��T*���4�w�_~������.��Cֽ���1�R�nndU�G�0�1'�i.x�Y�*��~._�hW=��.�=�P�ˢ�;���E��8ܑx�A6�V А�	��{x��4����>g4�	�]\.-�\{��Dɭ�
�=�D�;N(��ڞ���B=��+5�����ީ�_��*b���iG��Wl���D�z-2�d�>`H�$�#!)�!4vQQ����������oܘu0�p��B'�4���4+U��w?X��6�����|g~�|�����g	����w��kI�(��q��i%�b���D��q��O5�U�%��0%��Xqu���-زq�61����O5-�fi����k��'�P��g'�ce�׃.�S;eI3�MO�f�g�����n�i����p�SRmj%O-G4�������Zhc{�>j0���D��e�rѦ�v��9��Dp��
Mo��yO�WF��#6�j(Six[�����M��׼��$� �*{�UPI�l�@_lw��[�5\BD�8�A��h�֐@;un�~�.�C ��@(!.	�	E�.v��e.64W���.QQ�-��\�0�O�Ą��|��Y�gFS�4���d_>��	�E���v�D���N�q�?k��ɱ��K�]O&6������D���<
�L�٣��.[�������c~À}U$���e�C��#�z�j�)�M� �6��~	|���'l}2^%v�zRҮ��Y��?9�#z�7^�P#r�J��ޯ_��:���s��?
�X�'�j�Z;`9����+���Tl�m��Nf�����ax��K���>��1�n�)���L�A-/���,��l��, Jf�z��{�"���jTe���fKZ�~��q�2�_i���R��}�4�'����"PPX}�O*4��x���T���H���DnF���~'n�B���A���� F�e����C�	Ա�6���
�~>���rF�٧P'Hמh�qs��W1*����[�������w�0�}N؟�C�|{ҥ�ŏ�[Y�[���gz%U�꥘��z�$�T�f�:�ɗF%8�cVɔ���`y��ٱG�[�{CkUش��'���ɟ{�1'��mJ1��9aͪ��B�Ͱ�"M��zI��4�Ų�v5�+}>�`X��d��M���8W^49b�Ӫ���p��Z����U��ۣ�5�Ϋ~��g{$����'s�S��
�r�ʵ����1��})�K�K���Ʈ �Q�ROX$��ʿgC6��ٶ��i�3�l��O��7���=X0jQ_Ѡ�����MUx6�����|���X&^H́7�
�L��D�Mr���V[�QX��
b7�5.df�kU����M�S?�X�'�G�t旲J���gR�3�>WO1�Q�szȘ��u��-�J?�ke�)��?ԗé�?3:��IIQYNwH�H����������������U#�5�K���]h>���#<i�Y�"�S�d�5�,����7:��AF��ӓ�^�����p�m���fYj���Kϣ�+�C5>��jW��պb%��/EOic�.�R�B[A5���3���
3b����ձgKB��r!G�����<u���.�]I���W���jE�k�._X�`�3�H���IL�B��b.��*�B��A�O1ș��~�vc��p�̏�-l�$�Ke�e_�jR�#Y��\l槬H�4�צ|�#��[#5��Q������4�&��(f-�\d;WੌY�Q�Q<n��Mml�+)���p��u�|h�[٫A�x�@��DٿX2''��ӓ�f2���_N-��`㕟��*��[,���=9h��C��J���F��:P0�M�����������`�@B�S��@}ųFܗ@�JX��o����%T�%
�8nI����.�J�9O���&��cփ[�;g��\�7�au�����&kb��U�����`���D�&�P|�NL��Р��C,���e]�*���.�5[������v
���}���lmR�͛vR�X�"V���u�;�IB��/%<���.�_O�(
w=�LyU���Ù�\<W[�1�	���&���#�&E���ĉ���N�s2��-�1Q�`�Y� ����pi�V�G
�z����r�mte;��вԍ@���V��SUwᏦn+��s�{q$w~�o
���u��A2��֧��Y�^Н��)�"W�6M���W3�X�u�i`����Ŕ�%�����\qlX��P���YhFV[:�s4��.� o�nv'��iy'�8��Np����ɧ�<�����<� ���w#$Ď���D�y��+�+�["�8<�>b*ğ��UΜϟ��(���2
��i���bwr
�m`���c�}�2��
2����@銕:m��C,�g3�{{u�����q,1t������I��"�h7��̺���_Q*��6��c*g�oȵ��i�(�V���۵�A�gx<K|����ܶq����N�������\�ӭ��W~P���2b�A�Щ���b��ѷ�&��(�Ri���5j'뻝�����JT�z#�, ����;
��p4Փ�r�|5�7� ")�C��K�H�PNt�l슦�z�
hB�����o
Ym ��V��]�^�x��_��l��&�x&E�l�j�$����{��k��G���z��������%�\&�T����;j���������?6����fRN�Q��S1G�1oq"�ĲX;	a��_(2�Vd�<ۍ�Ze�?A�}�\7�}��lH�iG����QD��X�yFG�K�ǀB ��BЗ�����S���h�WK�_t �C��!���G�E��ޖJ�O��o{�������z^�Kc�4"KfI����������H!��b�m��ub@�jh�&��Y�ڕ���-�����{�޸�]{$�H�@��`<�
��T��͌|ۘ�}�i������]�q�R��p������F��\C�����LB�ȚܔZ"�B�#�ƃ^�Iܨ*/��SE���r$g��f�M��F�mMD0y9��$�݁�OJw�� �#���*��.������
�՚5d�;w�I�7| ���`qj�$�܌q[�%��Bt�?��*,�"a<��^����5g������<�ug%r]
����Ҧ���z�l�nl���Z�Ը35���Xl�����[.i왙�f3�� ��˾9u���>(3���1�ٍT(Tء�T�s���oSB�~�ӊ����Ѥ]��΍�=,//���3+�F3��9o6-���w�{�����]/��K2�����܇L�7�A	�x��I�K%ץ�1\]�D�H�&-��*����O0+nl�"4����1f"2ۦ׳3˵������M����[ٯ[���_�+����]}�B�y��!x�c :����
6���-9��aY<GR!*2��q���e�E��Vc�Q^9�?B��w�4��mȥ���!�tu�<�U�[��Wײ�_]Ӆn#x���0:Kã�r��i���[��+��癔�0�=HUs�E�	QP�ӹ��E(���^d��D�iU����k�{�� {�?i�|ÊP���a��yZa��4)�#m2˱��ƉMk.���־�Z�<N�{LꞱ/��,/����X]�[�,��/�6`���'C�|al�_��=������D���@;��C��i�!´s���t@�����mJJ.�׼�bz%^�YNg�t�����9#H��G��(�)��(y�S�ӿ;o�yQ�[ Kba�*�8���5�����\����O�3,�kP�-F���1v����ܕ��4��K�=����$���iNK����+%v���n4���+۔䜄������f�{~��J�!I>��d�=�M��'�^�e�yx�Nu����<���1�_C�����}��956**�����~{g���v�m�¨��Ն`��ZO���ىD"������
~Mq�n�q޳�o�`
��S܂�'�->�y�%�L��_5�3�����>##C�)��R�Ѳ�>:&f4��Cِ�"�&�z���b�pggg>Hc0��ʋ/X?���6�����_i���������0��0�p%�w �v���C.����?<�������W����ꥩi���x.~��]���3���\�-����F�U��X0��^W����r]P���G.<S��ݙ(нqd�PO�K���"�"��+gv�����w1		0���D
�f��.IvEf�$��#��{�������J��ûFϟ�W^dLv�q5�QRZ*�
��Y����7��,0bk�0Le��FGg��)�0�lwr��v���.�wFrE�E�M� ��0�G��;���y[��1���+�c��+�44\��p�h�3[A��aj_�z�V���Bz��57��~�6�c�	�>55o߿�Hy��B�"���K�[\6�i/�������`'��U��E� �?�Q��ty�4W����{,R��'�ˢxg ����{���	�JJ��������V�����bӀ;�_C%����rT��#ݾY(e�؎A^ߍH�B�|
��[4���A�R^\5H����!�s�=�̔�����w3��W�.%��OY<���6LNA��u�,!�[p-���?ن�U�t�D�w|g���Or�[���ڲU�^�N+h8���hg�/��<a�ׯ�������E��[m�.�?	��A�� ��ۈ��y��?9麿!g�EWR�f�c�	X<)Ĭ-��t�h���V����rz����0�/Lth	Wwo��A1>��s�䉡�&&�������-)��0N%=�|o}�Ts��{[�H7�)����o"R꯲>���Z���Cn���y���z-�DEG�B��^}#���H�,A��Yv�;�ۤ�
ȕ�A��̕�HM��
��ͤ��O�A�
\�n7��H
����$u��K���$a0o��c���c��U/�8�c ����[��H"�ߘ.{��N�Ĝ��J�e��ћX|b�}g2��:�_�tZ����7�}r�2�C�~v7o��Y�����	��s���Ň�zol�,�Z�q}RȆ�5��W�/ffd:7t����l	���kx�Myw�N�&�w�����I�_A�\����a�V�S�߯)���%Z~kM�5��p6�6CF��ޕ���.��//+��ɑ�m���)�˫Y[#����k� ����c{w7�|HF#����BX>���A2���5'Ǉщ�}eu�
��y8� ���, �?k)(|������r����505�p��Z�b��}8$!�k��1yR ���z�� � ��^5g��V��/�eZ����' ����]]��	I�l��81lׯX5����@s�����,ׯ@|����'?܂.� ���C";���7��b�D��������A���e��6X�<������~'��g[k��ش8�r<������Vz�-O�dhg�����r�30�0Ը�?3H������}�z,��pRDꐈ
�!{S�<^��'N!�ۃ�8� #/�F��F �X桦��Pڋ/�ZZ�iоT���:��`�����ɏTփyz
rr��1����5q#�- �d9���v� �^=C�er$w�_%�ڈ҇ư�1)�,�D��n�~�l�p۬Z���E�"�+e?�̷J F̊����Qں(X�S,���g3kyy��^�_f�ANEe�h�V�^�v��h���}���5L!1��d��I]A�W��^r�* "����G���}�x �]7;�]����b���ؾ�X΁~�� ��g���Y��ׯ�h�J�D�������9���	o�a1�?�����A�o� [��E� �w�c�Q��{?���sm��/�YV������XE -Z��8�@r���l��V�ENN���Q#�|��*���ÂժirsssB�P��,V��Q+�{��\�	���l�qq)��[��9ޟ�/Ԙ��L`i_���;ޏ)dcg�R >�0�z�6� A��P�O~<ow(����U�D�0bJ�ޖ�`jH�����ףȘ�lŞ�+���2~�zlp5���	�Z�0eK�z/0f֝r���|������@�^��߼�]�_�K�H<F��nJ���纒s�P����%(� ;*���5��{����3��i�ͽ�=\����ht��v�F��|�{�,��z�������%������#KK��W%	$D��i����ז��,�s�:�mJ�����c��C��z׏(�<�����#D��Bo�<8����;Z����&�R���֎p.�W>d�KF��t >��zf�*#0��G�T$� l�~y{{d��v�oi ��5Rj���G ������c���aQ.�������(�$�$-��H���>hdYn����sT��l��dm��j'\'i 6�ع�U���ө��7i�L��3/�0����j4Nn�w����.@��0�ȩ����
�a#����˭�Z�r��O�����rG�u���iw)Rk�3,!���a <�)i]q�-�+�������r,͸ދ�g<�Iq+s$C��i4�ߟ�h_#��g��t���!��l���@�R�i�P��K@�Y:�U���Υsa)i���XB��77��}}�_~v��{��\�9gf�����ة����힄��㽒c���<}Za���+u=k^H@ ,����L�ww�u��h�=PkdL
�[5j�����0iTE"1e���CzI��� ��������)�4����;��x��h���fhm]1�Dշ%���i�1�z9kk�4������?%Zɱ��Q�6��g������x�#J��Q]�z���r'E�WLO0?)�w��Y%��2K�,HB��\�4Da0[7[ί$�DGG#7��f�w������_�Խ��b��࿷�3���	0Μ���oP'	;�U��ăΊs��Q;fq
���+����^���n��Ӝ٫歟��d�D�:[˂�X��o�����Y�P����	֮{�zc��U��� z���"�]ޞz|`N'�%��������Kos�z��kKat����q�����#��3�N���1��#ݜ��7�>{�1aL�7n�|>豴 ?��bhC�\YuJ��&9|�����m�zC	:Q��h,�ڧH@D�m'>�)5�#	\�04,�}o�-��������[�33���1s㞫b4�� FDW��}F*-kg��p(��ID����<��-3��V����{�m�Zl�#f���f�}C�v�P]G���K ���\�ǖ���3�+..U)/&	/ہ�$��4D�������\�:�#/e�m��ҷr`d�ʔ%r�F�B#hK�����Y�}�8���;�ش�2��p�Q���������A]� �p�.װ�vGeJ2���i+x�U��SZ��F�jt�Z*ae�׋��`n|o,��S��(%Y�����A$�ra�y(c�Ĕ"����}vM�����#�mm.��(C����	��Ŕ�Ə�$U�uYRJF
�5Z���=�A��w@<��
�`�<)��<ĘGg�C����V����}:[��6PSS�V�T�S���7��"��3�����mqyy�ؤ��ֲva�d�n�՞��!���e;z��ׂ�.:�+�s�I�2���eѴ�
W;�E�o���L�_~��*r,ߙ�	��]I¼�0�f��~�$R�SY�-Z���&�"x<\i�֛��0Mf��&��P�����n�9Z�
�1�@��QQdk�U^^�>�� �d�Z��8�?l���
2���]r��nn��եN
��O��G���a�_��'b��Π{s���8�P9�ta��i�DQ�E���/��y��uy$b�X��8p]eX��|`����\*&�3�ܖ�Q^M�vg,7Y�p��QA�Q�^Ȑ�_ߐ[Q	�{�0L�?$Bُ���ގ1u�ӹ�e:�7b��Ɨ������)흩}��nP�.�'���rd�b+�o'�r�"0��ZaU H��WX���D�����9p��^�^��T[�����HĔ?1�s�j�f�JW��򋺭���%��qI�h%Q���#��M��$��?�^6�j�,Q}U�9��t+Q�����$P1�ۜ;�;�Ő]}?s��O�UV����x�_���bg�m�w�#�s�����J��$���w�.\�r�֦qΛNu����(湥=&n��z����ꨞ�^�����d����Bb�O�^5�����}����{�.a�TV�cي+�����\7�'pڍ_\��N90���?�w�_翍��w&?��*��z=W�~�L�f�{YKS3a�q��'�GG�O��gp߀�/㜆��g���������9���x+�.�4)G�K&�z��b�A���$����x�4���D����7~KK֦ff�)d�$+��۶��{*


��4yUw�ڙ�$ZH�AZk�q�������.�7�#��`i�=:���q�c�]�K��W�T���ފ������,9g�w�g���y�q;��K��cȝ1�kso�؀���U��3e�c:g�f:c1Q�7�w�BF�&����������<�Tq�n���¥<����l6����jQ�B ���hhdo�����>;� l��T�Xd��m���k�hLv�d�s���W[�F�6]�����{Ƕ6sU�@�C�?��F�N�h����kL���&�O`q���{t��k>����U�5I�\��2��-p(C���Z�gנ�����ڜ``��g#��x�@3��UlհU}��Z+��ԂYt�(%��Q-+0Ԙ\Ԛ��V��㫊N���ߌ���xwN�^P�K2�����g4����C�$��5}�PhtAFƃ��׮���[���.�7���z���9���a򡆺�<��(�-o!���gYQi�SA�e\tI��q���� ��!���g�ZG���V��sS(�Ew�Ы�{��2����y���򋋻s��_�1�geee�@����J||�����Q���P���*��Ά��7J B
�C�G*0t�r�tS������ƽ<g�䟓�jM�7u���5z�����X�܊M�t�R�P����"�I����;�%(8Xع�Dw���B���X��+�184��O��*���%b\��A4�L�0�%�t63'a.����8�K%��ƿ���lsF1��(� �R���[�3ZzX�c��Lr����+η��~�9G�e&�Q%k����,a%O������տ�`���\�����}}��������,&�����Y�;��%��߾6�L�5k��5Z^X�W���@��<X��H|Τ[�{� ���J�LXWt鬝��#�Hn��{���/��8h�$	<��<7����͎��3� g(��41�趴��~j��M�2a���E���\�PA��ٮ��$�n�/��&<1}ڴ�#'Ɣ���3�tb�1�7o��<o�f������e
SM���̏~����H�������� Ԕ���1%S(,4�^ef�ۊk��A�/�x�
��q����3�����\�CSZ3��/t�z4��Z?����8��c��sk�NJ��kOGG��YYپ��Έx{A������rOr�'<�9��r�j��ovM�c����F p�!54����.p�&�?;r��?_+��$�䶓SS�=Օo�Y2��4;+��v�``�g�}�ll� ��(`������=qrZ���XQQP����R�yYY#YU���b�g^\Z�hY 3O�ɇ;�yg!�Q|�a1����m6�.9�_'��C
��걸a nL���m~�}�R�/V? $$�oH��@��#�1��������(+K>�P322�-9�|}��D���]�u�\h�^jjju���}��i�Z>�o�P�CdsP�
��|Z***$�.�3��S4�/�̸�I^~���:����ꊒ�}��g/ ��V"��ɞ����t;�KX��3��_=��^��Y�]���pxT�y
�Z�ݫ0���	C!5�������gd�;�q����M��R�r�7�&��ݫd�#Co�"����7�Q�ۍ�ʗDƯ����CWV��Y?O#��u�fkO��W����n��d>R ������Z��,�Ç�̓�
�6Nt,�ā}�:�sF=����e�,�6٪�cj�ι�=�{*f�ך�7�?AP <��V�\���9����X�%s%#�}����W�wy�Dp4觊G]�իtn��&������b���1��-��"V5�&pv��l�P���6�r�� ���9KH�;,��`�=������r��oO��yq��CMU�����6���в���%��2_9J���K����F��~�A a�2��>�I�G��G��s��B��m�V#����bn9�ua�~��&?���$��۱21	E���lk�$d�U�_:
ḣv��x���b���喳�(х.�Uh+�D�hz�o<�b�g � ���yc����[�b�2�O>��a�^__���a<�]�x��a>����|��?��&}����i���R�_7hY�1&��?�@���8^�[]A�x�����X�Evv���Oo�iv�P�Xr_{���K�+���K��Z�a�s�N1�P��;�M�3���v]�r=�}���*����3��u���߀���.]��nh�*	����}x`��]U��{�@�CUE g�e�2.K�� �~��9���4�����X��������,���c�_�����ME�"�#�A�讟S�[q?�{��㖗�V��n7T��2>�**�r,�!vvv^؍755�F311��׏�t����OӸ㔇�@�cp��s�
����*�`�0מ��>����Ci�c����H�d�RF����ş���݋�>�fn�Z�u�Gu��R/:WY���::��:�O��n������^ K�1�D����	R���R�M>޽۶žG�Լf!�er�P	;fEDD���/?��s���XvCJ�J˝�0<���jt,��o�G#2?r�jR�R�!p�_�v�@�4q���{�l�����K�]e����Zʚ�J,�0����>����0�^��1�<�	M?�>>ޛ���(q�m憬����q���w(F�ٹ�m���s],,-��J �� �!bz�D�c!۶�=��p��T�#�Hל�;�L�K�,?�L,&���A��ϟv������
ŝh+]�S+x7�U��2s's�������k�m/�C�iY*����֟�c�{1�$!Y����Yl���0��5��d�og����� �zř����W�"�P�l�ߏ���T.$��7ꗠ4Uh[;�N;����+%�tg��s^�5K/�_���DϞ�;�E��_���`H�h���Uuu�j��x��["�98������L�۠����O�C'�<�x&~�}����S ��g]�:�4CЫ�ߚ�m���+��\�u{]�������Ko(D�'�������1�!�5���TZN=�}��K�/ķ6�r�J�0��7�i�D��ت�=�������e_��7(��$�ZR�W��u���&(<�t|�z��`m�QV��_/�a�d�9#��tɋ�6��Ŷ�"�����iR<Iʌ��A��5�\�bҁ/��� ,��w��m��6����|�`=C	߾)@�K����I�\��J�^�7J��+�\�z�����Fd��S��~��/ᆊ*�~||E
�����3#qq�ٹ��qm)���O����:nW ��ӗ�A�|���{�Sx���Z�t]�
e�<�0�G�{R(��ϜI(��[���jTB�A�!O%3*&f֕Ik	[��l��/(Y�������G1yihj��s�4>���F�����5�ϥ6������Ľ�(������H̥��\ۀ�y�	��^���PJ��:7-��.æ��۰�N�
�P��XCZ�m9.��#�X0��Qm�u�d���D��PS3.��<����A���z�>���W.�JNl��J�Ґ�n��1V�&���^����������LG'���]Z�+@|-�5���FG����.q��L�u����uYwfn�s�e��#���&`~�{�ɢ�I_DDu���m$����EE.��ő�`�U������.k�G�����gDm���R���|§˶t���c~����N�ފ_�\2Ov���u�IPǘ��cs1�a�m��7���ޠ���x�Ժ�H?Ҝ�\=�ma��}�3:.΢ �3N�^\���0)�ۯ��V��Ýw�E�1�n��xxE�������GP�n��:>����)m�6�QM3�2o�b��Ś��o������af!9�����e� p�F���5$.�a�N3����c���<��ɓC��{�%���#�1�p�b��T�a��XD[��,�x��5�Jԏ�t)Z�'�'��ј�������F�PTl,�+�_qHCCc�=+[>4 �Ɏ_�b�Z��������l���|��U/ў����Ӂ61~͙��K*k}? ������|7�1�*RsOP�����m|���5��_�,�ju��8������b�a��Bn���mѨ/��=�6 ��?|�xF��^�.A�j��ՙ�vr^���X4��~u��V��7Ԝ+*�A)\�E�|��'�l�E�u�Z��*�ÿ��|^�,XD��촶�����ڱ�I�Rg��Z}Iy��}Z���\5�+Ub��D��z$ե'��ӡ�P�$��S,z�wV���By�e^�Q�N�U �lF*U���܎w���������p�=ru�˃9�4���ޛ�����8�O(���m��KM^�eJ��{�l9�m��ûq��$�z�$���zRl
��XX���n�+M�>j�v�5չ�׮\�D�5H��� �
-H�e�|��ł5d�B��6�ￂr$������ؖF�%Q����Y�0��d'�՛��N��y�{�k>sQR��1����UwO>E[i=|�N���P��I@�\o}X����7�t���J̕��C2��Z�5C��*'�O�eee"G;S�蹹9A\����!~Y:�Ҩ��ş��r�Q�~'Joi`dgr�υw汹��M������ ��?���	 �kB�6Xiܷu��a���3OOo�1�uŀKoc��w?;ڜ�i��������M>\�~��0�B�P	.��`�Ք�[,��4�@�i�(�kdh�(u�}�q���ӽ7��i��G\��C� �T}�U�][�h��4���QQ��ͭ�e�]%��k�C2�v�S�4׭!+x&�S\�@�s��ԯ�A5e�>�������Ju Q6C¢�K�»C �@Ã��x��&�&F��^�OtE�}��x�����=��?�M[厦MOf��וּ ���ck<�ا`��PYZZB��Z9e{��cwfh=G�`�����k/��,}t�?π��� ��]'���i2��.�j+���e��<�l�r1���n�Б6n�Ⱦdx�t�xҵ�BO��?�����o��\\�Um��E�/)�^�V�
XR�'GGF{./WTٍ���-y{�n1ݝg/���h֧��cvv�Nq���kp�^�cv��X�'�� �y�`�}?�V�b;k���Z':���Z�'b7�٧b�e���a�Ϊ��Μc#�����+*B�ٔt~��0�hm���B�-����CV�5ؒ���i��|�m��3{%�#�|P~P�~Go�~DDD�γ>�]3��c�z�����Ei��i#��Iė�������/č9xO'�E2����ѝb��a.�X����/M��=�;�e%5(m,�r�T�Bڧ�����܍5:8��GGG��؁YX��w��v����H���
 q���:�^�)b���,z�n�}kԚZ�ۣ����*��*�����x��nǳd6�,SJF^�j̎c|k�*[�����������O��T�(&�w���2�``(��w"lhU�E��#�ڰ9�Gt�t��g��-f�����B�m�b���&[;�X�G��mm�3^�$49 ~��C^}2#�h�o~u����әw��D�h���� `�5���>��%����W�o��eG�� g߾}�1�꼍u�$FEeA-F��!���&��< ��XCBU#.>�Z��j������p.շ��� "��>�)&�ﻏ6b���-�W�А!j���<�z�4XKĘG��RY���p�t�JS�8g�Ϟ%�d\�
�l+*�?�L������jx՟�u3k���ׅ��L�bao7��AC�Ǘ����;,d򑉷�`��}�.����@a$�+�&�@i��k�4)6�x���6�]p��U� £s�4Ź_�+����BF��!��&`7b8%�^;� �Qi�y%%���P�h`	�Y~^�c����8q�=���|9eeD�
��+�::9�簾'����!�D��Oz���,%a�ElA���jq7�go�߈�;������
��Z�R'^�����W�^�D�`G���?�H�X�/�k���,T�'���F��R�P���0o3�ۦCW}�.~(e=��D��4}��y~ԩ�%9X�4wuy���*���K/8�k�S;�M��@4z�#~|f$� xZ�xN�-�F~�n�P�S���f�ʭ�K�_%�b�Y�ؘ�8�acc���"5x;�?i��DI�(�ߌ�,9O�)gp��Q�7ܦ��m������;b�o!!iK��m��f��8`�n4���97oy���[p�n�~�O��O�/��*��}T~����e����O��&��X	1��r�~��g*�]P'��4�Q�U�_���u�6�9������z���щV�h2�Y ��A�<��_����ׯ_��g?]�V��Nv�Kv[���D��S�=��ڭ�~��A��9o��=ū��/�����C�v:�$�V��n\�u_��3p��
F�#���;-����Qv}��2ڼ�ή�E������k+����?o@Y+�B{w�2Z��po�S_&�����s���މ����vq]]���E�z�,o��a���RDD�%싩P(�h�^��#�����~��&�^�vc��~�X$'$���������L��*���J�zw��L05X�qo�b����F@�����R2�m̽}kp�o}�h	Bϟ/5<T����_m2�Y���i�ƽ�fл�6��\>��4�Е$�V�t���}C@@Ӹ-�Xt��eB������t�������`�[�5������X�Z:��.�#Z!%��!*��j(e��_��s|�4E,���̓����u�X�������'�,��P`��G�5�q]��v�p���h��Pih'@�L)�UUU���
��1@g��zr�k�	cl���c�Pgp<�9$EK��89ݰ.� p�<�JnPpp82G&�^d.ɉ�uI;;7W�cU�L,�{T����^�-~X��vZ�;*�m�c`j���X������*@������d��~�,1��旃:��G��@kUiїaV��M��E�xڪ^.~�������zΰ@�?5-�~~؍�S5~/�r��N�6@�d%��@�cq�E6��h�9+��~
���2���៉B��1<�T�#괪*��5�U�99����~�hF�8��Eѥ�����eJ�����,Y��(��^�}� ��nb@ðid��,3k���|3��_*�덙>�n:ևz7�%������5��E��~bjj꧝�PL�i5ߛ^�����G4A���*�F�.AAA�:�]�~ �#��+IJJ�:�$���q��ˣ�v	�`[ۏ �.\�k����рF�v��p��߯�{���-y}�����atR�����#��W�5�l�w�#=O)H}2D��g�n���&]L,�0_��
/�NH�䐵��T2���<�}t��O]�����;Tl��{��1e��a�:�{&V��|E�Tn�� ���#����=X�8X���2-���Й�2���U�����J�l�7�������5����j\�Z9�%��Yf ��ZC�hML����iS3��'��)B.-�_�����r
ҍ�</~ �q��g����B$w���&�����S��"�҆��8����;���*�P`D�8\�뱵D5�<�]��U��,���???�W����$�w�y�l	P��ր�Ϯ)�)",��·ՇY"��#_<	s짠͕��@/g9H���4��M$�ώ���w*{��� �>�q۱E
����c�|9p�,˨G�3;D���sY��W:+�-����UZt���L#����׹D����Ÿ��~+�S�ɾ[�wuw̯��y(?�z�©`a��q���{��$���J�A���� z��(ʶ��çO�}7�,!�Aع�~%���D�6����oC�k�B�[�h�������|�j�#R�H�D�|��!���ˌ9��\t��ِ��p��=ܿdܰ��1�72��O����"W��)%��l�5�o4�����{�9��
�Xϰ���H����-�=}�w�}�ۗ/�y4$8o�t�٥H�:�vA��)B���޶{^�	���|�AW/nDr��mQK����i,� ��)�#��i�~��ut�7����G`%��+�ak�P��y��W/9洴�pP��h����t�7��3W����%�ħStU�թф�7���*�K�kM�kb}���\�E��!�(���� ���Y��U�(dS���Ä�UZ2�s��s����[�2PH��M�vK��JD��(��ɟ;��J�kW�C�~*���1ş��EP���-�X�Y�)�C(Q�*���S����jjhd���>�`_��4ڏr|��[�=�+f�� ��������||�p����6\�j���lؤ·}���_��U+��v�mX$f頓��t�K�/S���<A{�0N#����yt&�wA�рqcw誳���r7O�v/i*6 v%~Ԙr7���
l`.���eg'�'Y�w��T��@c�W�b]��|=�>���: +G�(�|�r�3d#Y,���7$|7QP�:�����To��Xnt���q1
���1�BN��:�4��c����N��c��!�N;1��+�kK�@S�x�	����1��C�{Q����х��TŬ�<����Dj;��0�`������	�>�l�>ɖE���ܾgn;����bȟ$��>@���_��h&��J/�k���ߩ����-�E�zaº~�)����1v^�Bå��ah.��u�J�
�������(6��ł�Oo���Qq�	l��[K}@睻p�Fu��e����'a�ӈ����x�'����q�r���E�8"l�z��GJ1w�?RQGw�*���!�ZVld>�2���ph�����W�sJD����� $��"J�JZ��$\�r��w�U�e�&+Z��~��O����'�s�� ���(O���..��VL�kih�IH2xo|ߛg����ai���=O�i���`Wd�/�ǆ�KD�lOߍ�8~�4���5��O(���~��&WʘC)�{B��v�a��'ڥ@;3�C�O��w�}L�;:9o��31⩶fA�!��Q
�2K�.|�B�2Ԋ� Iu�Q�w�b�3w(7��i��R�g��ְ4S_�ؘ�iQ�P��5r�Q�^Hqڷ�sfD[��v�G1��<����m5�Q4�$!h�rp��hTu��Ǌ����*�?��M��x~q��l�g�Ib�?Eبs{���{l���t���ԛFC�@�K~������`Iw�<=DZ��|�^�������0
�V����E\�jjj̖��7o�a�j,X!cjk�8���E1>PR���t�$Z���w�Ξ���	XO
W�C�����-���%��Wd����m�^����Uz�4�hE�̩I������f��j �B�딠�7��x���#m=�ͦ�k�����!�]
����	�u$og<��Żt����G��b�����'���T����|{�3�e5����B�T�e]�8v4[���~�����"k�Ey�v5��z�i�x9����zš�JG�Jp�V6h�Z.l�L�3-T%����@�طT�������$oW���>UŊ+��-�*����܂��h�͛T9Y�+��Y��t,ߙ�'������|uF��v�m������rB�@�ʊ��dfa���RQ�1��2��"�������g^` ,q��$�]���������eeT�Р�p-�5A�i4
5��e��Z��o�3�j�J'}� Lɲk$�>HQQ=�����+k2�����V�^���D~�f'�cf�H�[�N���m�y��L���j�ԻV�E�G2-nw�n�`M���M���E�d���
�(�dLц�'���J.���6t�^��c�VЩ�J��4y[A���6^������I��z�$�W���`(ȫJ�R��^���B���F��c�ys�o��Jg?F*��0��?�~��N��C����w���F���F�N�ɢUNsJ��7ђ��&'�_�v���dgԏ�7��f��O0��u/:Oayй�����G�Mv|w��Vl4y���]ZY3�`1����{���u�2�[C����t�����%���<�=�OD�0-���Z��n���&m�m��"y?�G��O�xގ��b�7z�S�k��'>����ȝ;SL]���n��t�����1�5������f�+�FX��^���q��ѧ�0A�q݁X��p���`���*ѬH%1��f���R��y@�a��ٗي��欟��o�x�&�Œ���k�iД���0�@�P)/�qt:�4��!��ɯ?����-g��!<�C��Ŭi�#}�3g�P�r����*{��%��1�9y#ݷ<�s���C:"��$��Iņ<s�DWZ�w�\6�7j�Q�E�&M�5\"_O��Ú�dC���_����:�܇�[+�S��]�Ll/�$��39njj�%�7}���K�Po��__�<��2���{���}X�+k���n���*Ņ�p7���bu��M�mV.��,����u/{�㥊�B�ѓ#2e�
Lp]�_�)��>�k�*��縇�8nc�<Ǥ�n7�>����H� 5��mf�f�]S���=�>dc�����Wm��
��#G�d��ͷ]�PM�i�3+�N�O��W��8�Ǟ�#���=�~O�[ߟ_�<j]�=�z�����-�Dad�VƊo�W�l^�g�?�ua/��(_�hƳ�Y��Wb�FNn,���m����Fj��0�x��虧/W�xļR�qC����h��������8l�8�T������c^%I��s��c������.��K�q���ϫ���+A>�="���$�%�r���]�1߲��)�L����1���ҭ�Q�y^(hb����r��q_�q�|J��b��W\{Q�(>~�"�:܇2�.y%l)��,*_�[	<��AH�����ҕh��������Xw�<Y\�KI��#���=�9��g�V�_�y	Z+��e������Lr�'G�Ep�y�-^F)֫]ۇ��jY���va�ha�8���5t�����94��.|Ѿjfa�nCl1��8T�6 ��P�L�k�:n˭PqL)ds�ՐT�0V�2t~Hǉ��0mwu�S^z�|wF+֢���K���3T�z�D�1�%;<���$��pM��D��(�UFX�-G{�b�V���%�7���j�bX0�`Qn�l@����i�24�(�*���W�|�A�b�v��˫v���������qNξ�P���Vt�������]km]�n��Q�bIM���s{Ɓ�CA�6��B�G��Ӑ�����Wi�N�q&'��S~�s�2��w6��3��N؝6�+Z�:���oc��E-��Z)���4�E@�
�0Vߪ�5�Z�-�S���
=x;l����K[ ^�r���{��.qD���D��k��X��uU�3�bH5A tޕ7�w��¦#pʫW-�7�h���L�=�w`E�^�b���md*r��l���\��ә�[�cm��ϴ;_���eR���B K�+������%�]��+Ҟ����(Ĥ����s� ϞIn���c�����1�
�acm���?n��o0b��<*�g�ض��'����XyV+e^��9�|G���x+,�nP�S9��+0��?��fߝ�Yy9�����^A��v���������,��_����X?5�� Otn���It�H`K��s��Z�Qd)�J�1l-�vy�d�
soi_d`(�մ���u32�<��_��n���'9Ēn���{L�&Y� � 6����4,)�4��۲6`LP P�%ߞ��ʦ���,��%���q��T���3���/1�3��g.�s���5N�9�Ű�?���v��L�H�6N�ϭ����@;􍋏��W���Ћ~�x(D=ո��.{d�z�tYL�rC���G&�j�,ug
�0��q�����
־�;��<#;�X�V�D[�[��[46o<94��Y4�f���l@�H;��p���nrd{�c���l		Ef�#Op�GVsD���.WE����.�t�������Q��S�-��|_It#RE�#�n��bI��6�|�Yv6r�&�O5�Rh�i3��c{=$o�t��r7��.�w������Y��D7��l���WZ��E�.��� u�{�]̿%��q5]�Џ1N��$+9�f��?|�Y�'7DN2�gK>kXX����2V�q��/:ܜv-h��Kg���H1<�>A��Õ�1R�O���˚`�Yk<ᝦ|��\z���LA��x?r"��T�7��y2s�У��T�h?��EW�[��/ghX��!�閌��5J"��A�!�$#]:�r�0R+�bٻEt-��p�59F�}�Ϗ��������cco>k��R<O(,�o���ˑ(�X����l��.��>r̻d�@��i[%����)f��s���m���^n��j1��u���B�9Z����5u}��^��@fG��'�_�:u(2<�_w����G|�р�Z���w�`�1�#��j��b���əZ��C��Ag��O& �����p<���D@7j�)Ж5�r>��wf�ʵ>%	�b�jz��y�>�7e�c�@V��!��y|Vw�$0?�b���-��=�mbp���+r&?&����D���ʿ�X_T�;�!݈͜�U^A[/�W�����,Y�k��=ٮҌ�IYwc�v(��a�\���+
hFTi�)�;a4�X����O�Q�����"��ET�2�%��d�a� ���֪����r=�N�_
�3�_>�F��Mq������wy�ҡ�'�dBIӆ\��U��
���?q���u�R�5i��x�"�V�H+�
p����/�5�G�x�[L8���W����混\ʖC*�3�(�*�C�ve2�������뻜��,�tJ�3kWG��m�"��!�K����Y��1���9qSU��L��-��Is�1�K��~��]��p�Q&a��gБ�~��w�����)���W�J@71�x;� �RK�{rXѣ/��."F"�V�����GZ6f}����qK�����o|�:��ϼ�X��-��WۂzpE�w(����Ɣ��V�I��J�v�cg�M�ݎ���_<�C ��N��|ϋW!�[+�_X�+�����$!P�Y��%Ӄ�m���@Qek9u�z8>�'=|�BVK�c`c��������T?S�b	�������J?���D��G�qBK�n��gm�v~�f�g	"OT���5��g���v����d�DWf�f��F��d��8�_��|�r��L�;�B⁝_�WB�{��R��9��3�����~���ׅ��ۍ��,�yϫ�֣8�e�Ѣ�|����]d�n���_J��Ed�/���2���(��7K��e�BQ�W�A+�K�(�b�n��G�Y��)����������6��|E��
m�����|BJ#�.Y�௜������:{2���u'����t����74|E�GBM��v�wS�,}��yS�����m���QF
*R-|�?�SكS��۫��AĬ�7�A��˝��$xٲp����X�0��6D��y&K;��T�p��:�r7h=)Tv�?^�%��3˷Ž
JK�	���E�;u4wK\��d|�B���|���$9�-��{��ذ�g����Wc�#�ԇ���\;��y6?	����h���>�c���#�OJ�C��|9��;_IV�l�m��ܟ��S<p�c�ںz���G�5��p��A+���Zp:��o/ߙ���e�H�Դԙ�����n)"�i咯J��D����)��~~�W����8��.Q����0�Eo�׏=et�κ���q,$+�)v����ce�J9��/5����V.�0����wqR��%}�[NHɲM�_˾/&�ޢ�L<�z���G&
��Sg~9���P��X�H�K����M�R�GЕ�{�[|,^�obi@J���]{��t.�h|;2��~�F�9tnsIRuk�w5�	"���c���K�Ƚ*��{�}���uRM��CcxB~&}mJ{֔��'pS�z�b���l�O�Xa�Z��vp�纻l��m;���K�R�֠�h�_Ϝ+1���W������-~G'V}��Y��b�~/1���,�Gv�f��5��$�{�ə^�s��5�µ�b��G��+��A����D�R�W����=���������ݵ=�;S�/K��DpmM���7^�:���{~J��9 ���O�4�*����W�\փ7����SӹR�Ɂ&XcP@���UW6�� q-z�#��=?0���[Ra&?s��3Ȋ�4�����X�G�$���>�"�;Z�����8�\�h,WGWؔ�$}��mΑиy� �P�5n��]#;�I�L٫��=Zym/yc���h�ъ����_��A��W��Yu��/�uÔB�ʷHgX}�kE����,��v�fk,m����UʡnB���֭�}�=b\g2���!Js+H�vL;¤O��ZK�-��_#��g�?�DڏPS��D��<�>f���g��K��K����%�&�܎������2cj[��F���mأ[ }̢�DE8�>��/��2����K�o��;5ȅ��-/���֞\Gx��P)i��;�;��Bm��#Oz��<_&�^:c��#$�N�KZ��T�u%�n��^7��4�[Ib/�0J�?lg���YY�?��un%Z�"zN�y�*���gBFGy �x�8���y(�c�ԭ{]������$Ez���,-��2uO����Ԗ����z������ͭ�2�|f.�!�0��C�-�ŭ�OՖy7���Y�m	�47���s��~KL7J�xJmw|\��N=�������(��}��P� σ7;�^43*�j�Z�EHфzDXj�����h�\� ����hH`d�"�L�}'GIS1�
��~��+U'<�vz���K��h��?Sp��O;ig�B�&{�e�z"%5����b,T�!eny�B��n'�F�x�*�Dq�����Y�E� f�6�õ9>7c��8�
�7�IODUu�����x�^,�I�N�T����Sa0��E̛&��˩!�0�'T"��/��|�����2m�?SJ�z��XL̵4b�޶ݡ0�Z?�m�;!c|��eW����&۸*�t�|oo���c� w}�~�8����<��b�Ei�C܄IO�Dߔ�_w3����<�}�~� �L��3�qY+���TP]*?a��~�>S�냳)�A;��$�^H�v��>/�ft�bU �-��iWٽu��* ~GjRs�X����Ğ`�Ocv&�F|�N픵��ut_Hq���7���7MFoG��#���7�=��)F�}r�s�3+������Q����qU՗(���V��Π�DS�V��
��w�ė2(KQ��BY�6�e@�z�h`ۖ�����q(}����� �r�އGQ9"�
�������0� "�C"�C�
JJ��P�=��HK�Н�~P����?��\Gq�yv�u��ޱ���@w�O�0��!e�դ�x)�� �%����~G�m+SֿcD�)ǒVZvԔ�*t����Ė��h��%�z�\�gp�α�������L?©�5}~��~����Ǟ�f�)�L03aݗ-�n�':��"�"$����n���U��:y�5\��a<ܳ&�y=���t�c�ܮ��KJ)B�
l}����ģ��k�D{{s�h�?>��ͧN�h����/e�0�t�Wa�󔨟���,�,LU��`���"5�Wq��m5��v�]���Kh���r%U3�Т��6ZQ���x5�Ek��Q�<3S�e�\�A<���n*3�	�t	�t${N^)Z����K9[髠[|���SeN��+�N9�&��f�Cts������O��;r���z��pFL'55GY_y|���������2%e��ק$��33Un<]n�	{"%�$�x䢭�x�sr����²(q䬯���F�ECfD�wh�W��F��e+��馧���mp4�~X���2(��;��n��'���?���y黓�{�����9*ˏ���D�DD�?��~=y���ۮ�R7N�|�#���_[g�˧�t�>�m$'�h�u�*G�F��tZ�!*a}�.����N��sŀgޣ��s_%}|�t�Xӿ�ݩ��Ԓ}���(��b�#���k�b-lY���j]���{-��iO�$���'6���-��������ȕ7k�9��ST�6o�#^}�67�֪��	�QU�JZKE�N^̃�X��앖י$a>P`ZXT�=��E�!$*
��"��u[okk{�
�����O��|�Z﹞t��d_�9���������ʗ�d�	d�� O�RSM���<Gax��X��l���� ������)6�?!�����h�η3;�͆�<�g��8V��qV�*��n���R�^����OO�~�N�G���4識�	�����]p@C�4��>W�`���;g;'>�ꙑ�J�!RIv�rJ_�5߇,^��-�KEdk�ol��Ő�_na7��2?�w��"��gG1%%%��8�F���S+���ȣ��67��糐,Yʆ偗����#��E۪�;�g�T�
���4t]�jڵU'�Q^�T:y�Ŏ<�nw�ל��k1��%�1GA�=s��r|}O?n��C�����������E:H��RƊ9�EO|=龿�;^�:�o3����xW�,�\wg����t*��cU�!����r�;ꍯM1L�йp�d�X��ϞV��v}p�������$��3.r�,&�h�숖�ꋲ-��7��z_m2�1�p�e]#�y��Žm��P���[�����ѿ����H�n�@���[����U̐٬��2����M����~��]g��L��z�;��c�xZ�|��Bx���{����m�$F8'��"�a/���no���ew���C�����@��aə�H�=�����{O�vT:�dcg�K�i�$��z��qKJu��Q���)�@b�С�T��B�p�h%v��:e^o�zΛ�J��ի�g������99�����i5�����g3126�x���{8_p��8�:LG�^:�ly��ezBpo����z��Tf�2_� �}�rm�D~̩nS.��㣍�X�C��P�1��-Z�n�g��v�x��:.�|�bΔS��fOr/���SU�q�	�癤�Aq��2��j;�w֣���6:kI�3��1�8����ڶ0(bQ��4?_�j������B�?�GG7�bg����pw�t^"nV�1Gm�v6����i��W-p�:����UG��l�߫x/XK%����|�;}��Ā��iB��FP
I%�J�j��K����o��HZ���9�N��s�MJ�oX�'��^N%��52����ٟ>]y��5��ٳg�deU���P�J��e*1�󽳝I� �����}%�膙z��N3nͩ�vF1k�YE1��dnH�e���R��T�z��~�؁�����VlG��D����:���X��[�x���tFW�L�s�q�b��MwC���܂$��c=����W��������xQMc=_mix�:+.-6�m�߽���|_�f�-�Vz)))��ϒ.s�ƨN�(?�f��$����l��G�s.���p*dp������߿:r)|���Q�]"(4WUQ!ϭ<�0"S��.de9�O��up��V�$i~�H��xW�QL�~7BG�Y/���Տ����j?z�X+F~�����+��\c�'A9�A-�����5��pB�^�3[��p!\��R0$�|VVpe��
���)*OM_i�2W����8�&$̬˲xn��z�j���q-&뤊㐰�.v��k݈����{̓���;�B���;�~f�U���.]�R������⒒k�q.�S	���XM��@C�]dӆSf�ˉ���Z	OxE2�ߗQԽ:���x6��5\z[h'�j4_b{�.
�O��ʦBBXs�:+��>g��V�Z�ІN���H����zO��E  �
W�"̨!�I[�g�;}��1���������&(6�����t����Ԫֱ6�����i�Si��L|��U�9�
�z�06x�����!�e-�������#�l7͠��5`'�\���5�{Xoc��;N���W�i�SSщ�5�#I�p�_�Dn]��''�=/}Æ'���Q���M�X����r��D M�q)��,���������$���h��̿��+)(���w;��I�5G>IUԷ�*hI�_�G�j�:��MR:NTy |���f{�q���M��WMM��[_����<�<łh��ݪ4Bn��e�u>����	.]xC##3vv����H];�#+���`AAI���@GG�x��C������V��s*UP�II���Ϧ�)�S��[��54"���B����з�" �@׬e#�z\���Cm�*��߼�E�
@�"����"5es�g�!�zg�ݴI��Qzy�L�rv��͛*e`�NN�5��t&5X�k��̏�/��(��#�a�T:�a��2F#��V'����}������ԉ~� �ڝV��\a�S�� ��7��4���֚�(}��e�g~�JKKsVB���F*J�5\\\
����r��[B�{i�h�GN{ss���`�^�����(��껲�&�q���Ї''0ؙ�i(������Z�,���	n���8�,�|�ljr�\J����6�(����lj'�<|v������8���g�1ek����w��^h;��?>�EşS��aa��H]'H����g�J
��mJ�|�F)x��\�\s�=�T��"��>&�yn��s�����^=*�?�IFKkonkˮ�#�l-�|	�ϢUt*S�ߴ�N��zff���`�i��Y�MLL�i�E�Z����1}oK8�>_�3�:��g-�o2���µ�YK��,@�m���U'��C!���Ly�X�)H*.�P:�^���X͛�����C��tez�� ���.S���F�Ħ7)-�Om`�,�iM�I�c��d�l/e�T��G���$֟�n��7o
a�ast��IϞ�e솲_Co�p��qy@�ϫ���� Mpʔ�٥[���Yw�@̇t~P�����4E*~�����N�/{�+9�))��};�P�`0�DK'.0ޕ�.���q��)ڙ��Sf?�>Xמ�t�̃Q��l��Š�)@���m��5����U��Q��L��?B�.��r��Ȥ�.��\�%[sNŭ���=J&���
*z.pgCqqqӃ�U*n��v	t���s|�3�ɝ�d?�'�蘘�eW�I鸭�A�.
���`�fS�����D(��Jj�yp��6�?"]�e+���p=	�X�'�ɰ�)�٩|e<+y+�5��l ���m�U��[i\��V�DIu{���b�'��J��m�5���T����Л�q����έ�������>�G����6���8�h��"X���gɠ�]�Q<�>��٫���[=��{x]�P9֊Q�n�'�D�`sX��]�#��OS�2� &���	]	;i+q�L�N�Y�0�I�-8s{�f%�;�l-�gt=4d��:�����n#␕=��L�S�-_��݋�}��Ĕ;0�=��jA�MN}C�9U�#�th�(cy0�$,�}���eK`aӅdq ���d�B����_K��k;B�ef�+74)g=�S�H0W^�)����PϠs���,��W�AF�;f?{���2J@���r��{���g���od������ȶ����Bw�N��u��-��<���X6NH:�Ƣu����㊓*�cI,�I��F$+�_���L]�vH��˚w������R�G�JO��(�D;G' ���B�#t+L����ǏD$$��6_@�X;G���ܬ�CQ�y��F)���<���L��6g�1ܘ]-��&�_��`,�z�;V3\�Np]*� l|����I	 7M*2==�e.9���T�],����`�u=������D�=��w���:���R���u�Jlly�E>h?��&��o����y'�����X�Q^��7�v�^rY����xql�k���� ���QRA!�>�!�4�=�!(

��B�$+�סZR����e�*�k�
�������y[[����@�dC �2~�h_����	����e�&��P.l�h^ņ@���ii�j9���/Y�v��a�L@�2�����g-∁
	A��~�e������Nl>r{��)4bU<����Y���-͈&��a����#��]'�PS4�j�f�o�U�>��o��e�ͩ|5"!a��8���w��SOp�Ƃu߆BhF.��~��G���;Tj�������OxC��I~^^Hh�q��h>�V��ݦ��ϣ�Q�۷Š��s����G�gA(�L9���}��0e>�t� J�W<�TW���f���������@)�#��à��#�TPQ	i�����k���4���$��c�<��y�����H�e�QU;7����{����4h&��8�o���������z$0��F���~,�3�|>Z�?�c�w��Mff�s��uҺ�(\\�|0�$���X�X4]
������'�.�N뾡hYw�ﰥ����wƵBJv�����%^{i��O�����D���;�?~�o�v�A�J�a���m[�0�����n�.w��>�<��./����Yٗ�5�ώ��*֒��	U�xEH�t<�oM�[E����eF̹��
�M:m�$�nR3g��������9ם�O2�v�@��I�y���l�_��'#�A��&��A9j>E˺��K#�aoߺ7C5ej�;��?��V�4:������o�Q��"z�||@�� �`&��:�����	a�}��B<p�^������N��ged�EEEe����8w&<�O7��f;b���� %]Lc���puv�m�uo�(P�#�디�������c��^t��ӭ\Og:ߗ�WP8<UhgkUs�\�9�(D����/pT�����歳���Z��rX�����Ǩ�E~�����Jy���n�e�6�9���,x>V�$������/ĭ.��(_��X��%��p�[m�.�U�����c���ɐ^EFj�H�9�,�������//���:��(�0i%%%R჎���V%/l])�]�»ahr�f��f�z���A����2s �333+��������4⺜�(� � %������0l����C��T�n�Ny���0=��(�vg.���j/n����z�g�O�r��JHH�W�k�҅��bE+BG^
�ꯡn)R�6�O`���J*�:	�l�C)� ���>�~Ip�x�oݥ��f*�����N_�#������UH����d+]69b�7{�;�\����i�����B��j� ��I��K]3-��_���a�m="н��XHt����٫�9(��y�c"��r����P�'vQ���O�7�g~c��:W� ���Q��&�<�lh���3��@�#cG������O]�<,ii+|�������ի�1.w\�n�"(��ǹ%��ޝ
�]�^=�� ��͆�H8;;;�� P3��E�����Rn�̠5�;&���'�_�*:�}���~��Ya𘘒2�>F�?zA�x������(Y7\��}A kX��Y$4����3va��P��3�����D?ck�>_������, �O���������l&���lb�����6�	��?���'$$t�z��7��B�I�7����?g�`�v��ω���'���+�ڿL�O��w<z��UlUu�����&�ݻ ��!uEP��!�����"���KG��	@AG��v���!��v`�@W�����K ��=555��V��z}7��p�&�����ng���;�2�IL�խ��6٩�t�?�"6��>�e�)�\���kޯ�W��'����^I��~��Z%m�L,�5K3������W���x���Gh`7 �e �)��莾2#Ϊcp���fLh(�	+����d�p����֜��H%�N�y1@i��OC���\����{(d?����o߾�Jw\�p���`bb�����+J�?~�C�5E&^��]P��0�Gy-NDU:�g���ݲ�
����U�T$%�]fվ�������2�R���D��ds��e���A��o?�@��C������Sh��Flq�;���Y*��ۂ���VW� �I����4cFc�{��A��ցG��_�N4L�:��àZ�ȏ���Y�'r�h����\s4�V��?O���J�ҧ���> B*��c�A{O��H�Ha�*��T� +A��ai��(҇q2�͛�j"���|�N�2v��Ȩo�
4N��v�0��}�t��v���<M��o��u�_��G�c܎0�-�2C�Wy�gf����C?e��)gBȞ���峀ׅ&���E�9n@s�|]|λ�A��Y+��޽���-Y��+�������R�Ӝ�Ν��
�Ќ��؁��1{xV��!Tn/>�w��ֆ�
x���E��ԗM�m*�?�0n[
�2ƕ����H�D��Ѥd�9���c�h�Z/Vd+kQK]���L.��5�P��}�9pô�.�I��N��{�bon/��K���R�(fm����en5��!M���Y��$���PE�]�!�}�����:g2�455��@:�A��~�>H}Wl��T���ru�������B�	�`��:V��G|jS��c�@s=0�mk�q��2����Vk-bz}�0�o��$pQ�æe�+d.0/��w�Jcݓ$�嵜;!�ԙ]v��PQ��,�p�A�"��%iY��ǼO���:ϫ���?�o���?�N�Z����AiD:�cR�?}��9�������	�)d<6�4b6	��`��);۱A�>�^�ΔT_o�/PE����Ў�,%�g��N;�_�-<���k�(=g��4�Y�*Ğ?��͛N�ԄQ��{��/�J�&���ګ�?�F��-Gӿ�W�ɮ�ʟ�t�`m@����F�������2�33�����-��Ш(s8t��Kr�0�袬Ũ�H38��FZ; �Ƞ �	#�"S`8�w{�Z��s_$���`�J��)����G�Y������^a��S���RJJj����-'�δ��I�����3��MEG_��(wX̨���u�ɝ�1��(S����|�fN
�����MvҊ	�گ���58�i�<l���>�����i�9��/ t���c��|�r�s��K�!��d|jk�_� �g9��.����:;`N�TGc>�2��aa�	�ouuP`J��e�L��O�s������ϼ�g�8�v���.Jq��w�u���#��I����󞧷����Yj7C%�&y�I@�XRRו,��o�,UE�7�����޽{?]U���S�y�ڀv�_�D���c}���YYFF)�l�������y��h�k�N+�k��U��,���Z��Q����J�����+˥'a^����#%�v�Z0��B�.��B��1��3� (��ǁlLL]�g�i9�d@�����:��2��׀���X�q���M�$s�7���nb��T�%e�Mt`�d�9|0���8��<�hg��o6U��3wbJ_#B ~�Lo��a�1L�Z��B�_�f�&�G�4VH������[��������x�v�ܷ4b���9c �̫�o���՜c�\�ǹ���� UJV6k�z*ݝ;P}� �k�Sd{�$H)()��h<S'��0�m��N^T1��2M�}���cL�n�U̜��'I0 �CK�s�y�$�
~���t[V�}��"q�g`��(�щ�V��������%�t�C���B^���{#|w�e���p�M\/*l����)���£�1Vesw���`MH$5Km�M���y�.!�͞�7�0h	��ߺ����W�L�r���s�n�J������˓q�++�ec��R�vXǈ�?_��V*Э/��h���k������j2��=�Q�툶���B�O������m��^��k-y|1,�-E�QӼ��n�"�ksp�l%v�5q�Ń?[�T			PY[T3K�N�R������M2���-��>����l�K]	�UK�@e�(+>^dnn.e��Y�gI��^'0�J<ʬ�3�oM-2 0g���}������m;��)k�h���i�[�k�������kx�Mb��с�����d#�^3�6ו5T��=��H��5
�b5��+�{��;}�˯��֋���S�(����1Y?��UTټ�R�I�D�YX��0<q�q�\�n�|eS�Y��M?��^��0=<�E�,H4�bI��Yu�v���YF��(��r��o�/�(�Y:�=.�+d\�(Զ��.��X��C��^��Ք�>�9h�2ٮk���ߖa[�W�U�+��Qop��U�VT-s�2e��B�r�՜�=���&������n�O�Q{l��r��c+W��e�D.���z#�Z e�܈<D�
��J��2�A˾����-dgX�Un�:�3.��ܮ�t��!X�&�$>��<2b>��'`���ޘ�^r��$��+	Ə���ѣ���i4�,x�8%�))�1���n���P��G�?r�^�V�A_�iǂ���;�5�%lv����R���i��A�L���vV����xI��{��ݻ����-�5o|% e�Us�E'��>h�3�<���k�������w���|vnm�<QPN�B@Z�0y�?�
������5_��G/�t�@�DBe���0�{�q��M��xh1���9U$����6Oq]*mXUlH��i�}�a&;�@��#&o�8ם:o��w<��я߬��U�y�6UZ���=t��+����g�l[����I�2��u��3��}M��T��*�g�[�*�RD��i��V%cg�R-��/��z�QY���wA��}���Ơeh���5>%�E1��3m1R��h�> X��q�EP*d�V �!�n(�;�[���˗��8&;��^t��;�NP�)�� @4����񵚝�~��2
@���DF
��[��aa�tڛ�����T�<e?���\�)�ں"�&~��T�faׇ�bP�%&!��e;���B�;��A�YP�N`?B3��C��M��9T�����9X��
���hTSQ	�8PI���;О1�������m���@�4дR22*��/�z� �7��>�:�B�6���3qK��wZ�\��R,U��ٗkjB;�*����ʵ��j���
L�d�,xL/�SYo�o���E���^$���M��RoL��!o�R�6"̫_�>Ѹ����R���9��wo�v�0r�����(D"ev֤ФST��~���6t�locζ4Áy<Z*�b��J����Y��hO�he�A�29�22=��
�B#��CJ{8�\�l��p��T9}f�p�ט�Sx��;72�>��i�|��l`��鿦�����%��aHT:o(���Bu��kNe�cY19�22-9��{1�>�p�'t�ǘѪ7?/4:~�Lù���jO�Y�u� >��4A�p^���;:H�U,0鼥�4�*`���t)�P5�a�(s�b��YfT��P��٤�=績LN��25]G*�G�S�b2F؎�0*����_,���v�r|�����L��] ;,�D�<��/�y��k�9�
��q��/�9�\��=	b� ���K�Y�E��04Bn�kx���?F���O(,]p=��ۇ��.N�6
�*.2Q9��ʑ��T �A�.�p������=���U�g�� �P���k���C �鹹�O�c��	Pt�v^���NVU݁��f_c0=�����!L�)ɦ �4��	iU �&"�;��J@q&Lmu������R;�[K��(���S���`d��
 �z������a|��}��M�Ѝr9dԮ�E7&�r�#oc�bX���fYW�>�RE��x{cg"p.D�^DM��qM��E _�XF��["8Q��=&1MN����� @����o�/��A��=\��@� ;�K5�o�L��E_rTL*�#�o��T�*�q�[�`0�P:h�\��`�*�1;��j�Wm�����U(6@e�U�0��ZOmfDf��fgg������#�z/��c�V�].��	�҄	��h��lS]؄�b,�����9y�*����3�/%Ezf�h& 4�|���+�<�v��_K��� .'��v(�2�"2���eR@Ũ Ce��14�͢[���;]9գ0;'xho������:��������x(�4fUn���j����-Sggg(9T:Iի
�QeLmm-5��\p�����d�� M{���	b>��]�9��<Pu �T��ǥ�c��@Ȟ��A l��$��1Pq�M`|�I�����L�R�����к���F�U��Gt
*��:��Uĭ=�hk[J)+:�W���Ⴌ��v���#��f:���a�m��ƒ��.W��~�h8��j��%��y�J��[�P�\(k�p���]����K�h}�fC��2&e��QK��m
��A>Z��k^�`�M����C�'��Z�^�>BM[ۼ2����4�4q��О҂CyMM�������[�/3ݾ-Dx��'�a<P>r(��?~\s�P	(��B�CCCT˝�v���κi�$��F1ݙl�?��秪����"ch``$^�ZB`��
j��� #77`�Νn�4����~�?_��v����̵��� �==N�>��ֆ���&~Qߠ��`����+n�����"�W�� ���r��5*�eZkL�C��!�â0y��.�d|���h��R��Y�_������� �Q�V��J�qE�������Y�*��"��s�C'���~��U�H�C��*�W� n]eu�ǥ���hXI/(P� �}|n��dK_�r���u�sۋ�8��]�z��NE`#ж��L��j��������2���<=!65|��y��wd��PH�8<Tx	�څ�{���'x�6����}��!�×P^�tT�w��M��Ha�%+�פT?��搛i��6��7��_�1`0�j��x�����6_jλ�>?�#��k�(�/3��]��{���FO�Ӫ>Y��<��vc}G6l�G��0�J-#s���X��w��?�}�\C��iK��\L�Er���i�%e�>ǐ�2ұo0��_�S�̞t`��gA�J��H%n�E�TЁS�N4T�*��a�@�k Q�o��N��11��Y��񖆖�k�����AfS��iN󤜙!�xU��_�a^fІBf{(�x���F��5�����X�ɦ���x�u�E�69�&�KF�[���y�9]JS�u���1~r��1Ẇ,�v�I_n�jg�O?2~-��;�5���}����U�>i
�6�պb���D�;�z�UA�˹�sf��I���?&Z,�6����y�b�3?��[�~ H>yu�;�MI����y�(�}��Q�k����)�NI@���4�,��г�������<��s�I��p�x��ICp���>��������A��ar��c��C"�0FgA�ѕ�D=�*�/��H��>R-XL^;?���8�[q�'��R��~N��~$j��9�_6o��<�"���a+5V.���-?IB��_Ŵ��"z�=������t<��Ϙ����N]��(��V ok�/ū�"B�&����Z?�m��g�jJ ?��ǽ'@q�<��Hc�3��m+���y��fL�C[��rx�T�yʚ%z#Sz��3����1�^fp�o�=p(\xӐ@��G�Y�$n�!��`��9CF�u���~]* $mHtt�y�5���e���h1�f�\��l�8�v��ȹ����S��Y�p�}��KT��I��qDk��D�m4?bjا�<_��������ע�Q_G4Z��Q���s�[I��S|m嚆�>��w���Nk�J�[kf�]��D��PѸV߯��IL��P��D���QjҜ��z.�Vh��UuY�'��TB�hR;�ghC��E�젇dǻO W�Oga�z��F��lV(��c4DZnqM�:��oXD�~�ǒ��+��Ъ����y��*�W���GU��mu!Ӣ��]1�/���|�f��b���w�Y:qx7�+�NR����{
���LU�QZPO���f7���^	�y<[+O�b����zy7�z�|1�U6�bE'�G֜_V�/>r�����m��y�y���qc����L7�� ���j1T?���]�{�ȯޢ�1J�1W�� v�a^u2�^�Z�%}��k̖i:_��}ON<|���B�Z������8��z���c�:GQ�]�e�Nt���O:�
�Zk5�T���_�{�u����[��\�IةG?�b�4�	��δ082X��Թq�zn� �t�����^�ӂ]ب����=<��꣮��sng�|�(�D�'�Tb� QT�ۿ����\E}�U��S���,�� ������3=L$XP�<����'_����RĨ�t�Ǯ��*>��T���|]�[@��Bh���c_A>D}��]	�ˡ;�:D|a�(r��������|�G�A�h ������\*Z6�ˊfLJ�1�I$Uл�����+#]Ӡ��EK���'j$Ga0�7�Ȝ���+ оta8��l�fP��%�$�˃�ٳ�����zk��?gV��Q�zN��R�|x{�GS�)]J����@����[QI_���z�?���e�H�>7���!��k��(0�Bz�'��?-���/?,>[ܣP�>5�~楿��J }��-!,~�oϓ���NI�r��O}Y���aS���Yk�?m���O]0���g�����Z�&>`\�e4��C����W��~��<�w@���T��z�$y�G�⨵p�̀gj<��ǻ�B�l�Wg��5��&b03��jk��i���#��	>VS�'� �go����&vb�m�Wy� �C������WF���ܯ�h���QN�7����2�%�l���hМ&Q�,R�b���z��v�OL�G�vJE{O9�2&ND��j�"r3����~>��H���^{7�j���^���Pw����:HBП ����������8�`t�vA���/�Gw�B80#\�B�^p�3;u�[�ߨ͠#0�~H���z�Y�B��*l��h���$��Z'vdr�9NA��#�z��\q�$����a�p-��u�G:$���F�)���[�,�0��h�ӄ����ux%�+���w�k�A�OSXh`;�eq|��/���c#q�������W�g�d�S;���3��i8�.��n��jY�}b�)B�b��Ӿ�U����ζ�"��4�7�_�eIO+���E|
<d����לG�EO��5�#�����ݖ�^p�}e@��Qc�
>�;q������ω�tI����D��xi|�Wʀ`D�ԎA:���?F�fi�|d�}O�&4}�<u5�ͯ���� �S@m�R�Z������K�_~ =�(���4�J&x�1�Cs���"O�n޼s��HPr���1��p:��t��6/8k��b��/9~�l:�D���k؋;��7FPK�#��wB�T�p�3�nn����`��%�e�sLa'�8�Ϝ�`�+��b�r���4�A�If������[���,B������ݡh�է*£���ܦ��ϖӕ�����>;�u&=��ԙ����D%���M�v���o���G������_8҅��y&�}����-/���؇�O��MZ�F?�dk-;c
�_��.S{�|���=?�
5�Dǫ���u|v����v��(ce���p���0�/��a?JL�����J�6e,�<f��Ӛ�nT�O�x�{5�6~.-����o��d���B����4=(w7ۍb�-
�*E?�Y��|O0���V�+t���*1!��]�O
]�ʈދ�)��aޙ�V�]Jo��z�����75_���l��}�3�N�D"�Wv>_��0&�B�P6�g�����<90$�%�2D�R
�5!/p�H^
�3����|�S�����3����LMer�	�q�k�_�]Q~�2۩1�����k�9�g00��eb�g��l+ѧX��_�MBmt�AT�힏G�.�K����?V�n9>:3s���^cV.�禾8�w���>:zo��#�i�����0�3����_��H���U�t�9�����['>G�\���Ύ����K�{鳋x��.[�GnܦV��ic7�Q����3h�+oB�H��t |�m	>%j<�v�k�ve���x�[�������|ܲ�n}��-��5#U�~�K5C!��9�ش9����;�y�=z����L�u좍SAQ�--�EA�Q���0�J�?n�u��9��Ao`t4=�3%�q�8�%j�@�x$�*�g]i-ͭxZ��������pƩ����������"�݌���&5Ra�dN�[B����Fu�I�o��]R���VfX,̸z�Oji��oڭ�h�-r��|��"�s�����}�E����B��~4��3EcϽ�s_��\���{
ҚB�W�D����ϴ
�/
y2x�IΧG�K��j�3��Jta�Q�^M3�6�u���q�("��P�n�����-M5�%�6�˷�&?韙�ĽҞ�|�;��ׯ�5T����2�u�P��ݷ��Ԯ=�t[����X��V��_o�� _.ճI_w�^��Y=M�PU�e��������QHu�Px�>BQ-t0�"�����9rYZw�4��oThWI��ʼO�Bg~9O�77��n8暵~>_��L���nf}��SQ���^UXK�z��κ������{�dɦ�;Qj�	��m�F�C{U�~J�/m������IEtl���3����6�k�/7(�����Q-q�i���TZW+e��"Km|�]�΅�窅[�߭�c�x����=ףlvn�Ĝ��+=rc]�Lea���6F�g"'���/���
U�o�V���ی�g��z8�RN�v�`*�A.�,��j[L^�͔Xg_''L��xmv�i;Ayb�α��CѦ���q�[
&�żQ���8n�pt/��[��o���I�؁������w�����/���Q���1e�]=z��D��:�#������5��j���~\W<j#"���4!�_$�����[B?�{�c����'�y�V�<h�µ?Ͻ�����Ҽ�	���G�<�;r�q��7��������y/�<�>+�wm�R�-��F{<��u���$ò�e(���Vvu��� �v>�z��Οq��� �}빷�	$��DsR]�5�kb�y ���w��$w���,\]�d���ov�e;a7I%n�,�����2�Eƴ��x���	J.Ҏ 7�Rv&e�	��V�����G�S�ۺ�j�� !��,�xg�?�� �<1�����FFTM���褍�h���?|�����a��.�%�ݕ�F�M�\�R�c��h�����}1v��͌v%{��9n�E�!�͑���F1O�b=�_�E���˻݂^mb���߭psY-�%�pVAF�n�}վ?t���кGuv����9n�gr��e���<�Ke�M�g�(�<o�uվ�e�d1�FU�F�w�+���#k��#�cx�c�O�vo�ޯg����w �R�FD+~��/��{�	4�Kr��:�=��8�Y�s�gB��5�3��EO�Uj�},o^:c�{����N�$���k~&����xDA�'�Fn����M��S#�����Ky�#��V?N�+�B[Ԏ����"rt�`ZB׶�Ү<H4*�!���.�p�i��V.��l����T��g:48�~�2d�K��%o8�2���;qDe�ly��3������g�6�����JK�2w;7�D2P��Z��c����v��w�����D#���8�`=y@7�66�8��5$HN��!rA������]�`�`�%���73| �*n���@Ӭˤ��Ye��.7��?����h�1�����`�>�h��ے�Ͻ��K>K�<#�=N�C���O�a�J��[&f��(��,�ן*���2ɚp%I��1n�P{��6�U7;��R��.�}���d�?��7~�x�#P8�q�м`goY��~g��y�(��.���:�k�d�%���:X� �7�t�ZO&�)�'��/׽8r�8��t���6G�7�`���Xx�}NQ�,;X��!���lg���8�������٣����������S��4[��Qr��nK}��_3ދ��t�P���y���RΣ�#hr"8���]�������wul�>�4�f��.y�X��} ��{XRY��+�\�g�RY�Ԗ�a���Vr���	0<_W�]�ʒO��`ҩp��{�l��z�����llP��SR
���$�S?��W�w�����_��k�f���������Y��FܳepZ��AK�B}�5��t�YCN��%+�ym0�wq�m�*rnntWXXNrV�r�y���gI.nK)�U���d�,��
+m�z��=�GYH.	w��,X�S��$H3}�i݊�l���a
������Yƀ� {_�j�I���&��X�Y��x�����C��t�
)e�sc������խ��O�i<���	2���B��}��;7{�Q�6����v��څ��X��p�O��eGK�8R�<@��ѕXҙ�x�\�5���F��M}z�hƊ��-Yy�;=��TT<b���ե����j+��w\Qb� ̪� �=�7�w��6O}��G�]�3��}`a��$��`���,.tz������jֹ9߃zʼ6�ny��-���(ZSÅ��|��t��Ҧ#]����u{��l��5R#��7�3�7_���֭G<������Q9�n�-�V�b��)6�(҆��E|�|�^����붠rO���D櫻��7T*di:��M����,�����ſ��z�
(�x�AcK櫢�	��屟n~S>�j�7����cO�s㴶 ����Hi���v4O�;����[Y��`�f�-���6v��mvqjЇ�]��N�P�
� Ɵъҡ.�ع�d�dS8�'�g�#n��ir���h"�c�Y訲z�O�崁�ŀ���x�B]�������8\Y�"�:n[aa�mr�·���2~M��z(��ad�-���Ɠ��K��>2���������@Muk�Q���"M@DD���H��.�D���+��ދT� �t��Ѓ 5t����+��L�q���Ե����Dq���w�����f�͗���ML�L���� �b6_�}r)��ܼ�$i���Z�`{�&�>�2���V6��a*1mX�������-��V����}}9Rk�c ���~�M&���>@D`^�����S% _�����۾D�@g˿���6��`��o�^nn��m�<,Z��֧�fl�Qyfl���_+ALfj�6AɾP��-@� %�Vv�r�jv�]�0����Oh;~2�w�K�������uT�Y��6��}��qz�3X"
̼�_��+������<��k)�.׍�[߉��31�49[x-�����z@��%Ǜ3O,����>���c����n̾�)�e9R����l���1�"��u��ý ����,}����8������~��~dyv�ϢH���0�i@z/.0\��`/�t��WK�/�ڃFSd]� ��=?/��j��)'�J"������|4�1G N�1�8sȎd�������0����֤Sf[������,�bF>P�Q�m�t���E�_���1M��"@N权7�S��SR��Wm�ͭ����¯E�*����6;!a�w �����RF�Vğ]Za�
�&Eb]�Xaez��P��h����b�f���Y�����\y!���RU����R���D��n��d�OI�4��ծ�5ԍL���O7��8��nVy�=TI.�������O������)$����>	bylK�`}b�ȶ1k�#Y����	�>�Gg�n)���
���[?B�d��9������DgZ���D��?X(3�j����8��D��r���ݯ���LrpxU����!q��	b7�?��]jϠ]��V����E��G�~����˲D��JA��O����8��4GJx�_��V1F���[f��A���k[F� 	�G_4�S�--�.���+O����ٴ�S~g�%�Cς����@�����Y�����M�1�%F3���M<��W+DP%Z�����m���G"
&Dg��E��"���<��/˄sI�w�<�Iv!�?8���Oc�r5p$P9�겙�u(Тq�P��\N_���cd_p��:��:ъ�ݳ��;�r����8�s�Z�����R0�۝(W�������%k#������x�Ji}������Yb�x�+����3门5���o�j5���{�F�ub���A��V(����g���T��yfq����tt��^�A��#l����~�����z���Ϭ9	�n��
�"t���Qx�{ߣ����l��m��H=�w�#9z�����C�wD�)�|����ʼ�;��_�����1���Y��I�m�9$��|뾓׮olp����f��X �@r6�nI>w��¥*9o2�|����SN���jE���n�c-t�gX� ��F�l�1�o�i��6�u��6�m*�.��� ��"���ٹm������g���෈�<�k�ȝ7��P���Nz^�2�0(Ϙ�z�/�����ḅ�#pbӺ����/Ï�h$��>Nu�O��*���d��K�$�uüp��S�3;gm�-5S%��{;��G��䊱q�,%ƺQ,l�^��ϙ��\�f�~����e�q&����j{������zM](*�!AD��k�@e]����]�Ѿ�׶��?�ߘp�9#[�C�]��.-iSd��}�T�s���9���o�fFeD��Z�V	������oǕQڙ=����q�o�����<�	1ŐI�d/�VP��jS�Wո�r�F%l��z��/�%,�w�c�Ր�N��ON�pO���>���t5I�ɵ� 6�W�J`��6��]I���3�5�����-�צ�XA����2���?H§�����?r�]���j�@皘/��F��9]�]/�)c��'E�e޳,�\��`! ��J��x���ڸO���N_]��W=�8�S�.
�BT�\����<�������W�d�^~녺ףGWՔ1�w!n��$�aP��'yT���;$l��)g+mF����;sy�Dl���r�o*���uA�;ux��(�w���A�����"@a���	0ϭ������ ��e������g4�L� sTR�A|�	P�V�J[bzL����{�5+LzF�~�]�!�<N�I4T�'��l_v��	�;w�����%J}͌O�tܦ��w �� ?��+9gEe�@�A#wq���3�%
 zG�0C:���L�ē�|��+'Zl�KEتMV'��B����1Q�?P̯=�^�R<��V�>	��	��\��ܿ��8���"�vy���� ��Xw�#FT�J�?Ȅk߁55�J���r6h��Ђ��<��_�L_M��Q7Q���]�4��I]����6G
��!�%�N�0�ĩ�|��.����3��E�e
�`�R��31?��P0� �mAP�t��	+oA���I�mQJ&�����^uf�Y<����C�.. ,GW,Ӷ���-a���?��n�Q��]�buS��c��\�N]���1��0-����}�-gD]��4^��=�BV�uR�C��u��'؜\��z��YC�F~�K
0�d���X�6�67-��D9v�`8�<�k�KF�Z�{�7H1��k��ű�#�Ό=.�.!�$L�����'�:����ME�Q����ɲ�낕"���/��FD���.�(�1�V/1PFU�ץ��z��'�2(�`��MY㎝WG�OO�ț�1%��V�*�
��;V������fA�TP�$ى6ޙf ��`5ۄ��(��k�җ�9:� �/M���:=?J���ʵ!���B.�S��b/��f8� S؏Dw�pIW���?���7�sf"ց�`��`�\~����?c�ھ�Z�� ��P�r[Ɠ0G��M/�|��.�LY����=r��~���B�jN��*��A1RDN���*!h��&�`U�w�Km��& �&����1�D�+�V��/�X��NLg�r��֮�����Փ�͘���.
#����w`(� !�#��h)!�u>��&%�CZ'�<�Zk �Kr���It���C��h���N����eމl�&¡7�)V�n2�\D x7�41�`� �
MӀ����T��q�m��Aݐ��g`P��l�˺���}u�������U��'je�/L�]�p#I��͛el�=��hB4eY��[Vji��7�(S�%Ǻ�y!��U��,&�ƚ��|��@����[�������	���E�G��!Y�唇@��|T�>@k�L�z}3����aT�F���$��!�DP3���<q�^���.�oߕ�١��%w2�����z]*��3^��jw͞��2����=��N���h}X� ^�T�_��Yk�<��V~�bt=B����G����.a�Q���a�nģ��IH�.K��w�Y���s����E;�MEO�x���M��e[�R�>wc7��� g��&�����$8&*h,��ZoՎn".���m>�v�����Ug0��VK�nd�A��B��onv����-��sL�y�����η�
$C���C)F��W6�֕^����㱪�x�`�@F�m1���c��V6Ѭ�6||�}ϱ�K[Q�Ǿ�7����G�A{'��ktCf��{��� %���גվ��6�/H«P�3�����f�������79�@D��A̯*�_����ei`~c+���9���}�_2��u���˯~�IdÀj��טq���Z7����r=�[O���@Vht�u����&�8,���ϻ����C�m��Q_����0�3e��ru���+�~��P	y���E�i����l?�.�+e��g�Pa��v��j����2�Z�>`ҽa�hFJ�U�=��vР��K`�1I�48���8��v[ru�хL]�>�/��I�c9Z�`>r�j� �re������!��~��Є�09@��uC�a h��r�3�MgC�P0rE�r�H3t�ָEVT�vP���;fB�������Y����{|��z�u溪MHK費q�d�p.i������ʥ`��q1?b�*<��Z��o�����z��M��A�2uaJ�O�;�==�*�'��Ӭ��5��aKKߥ�ї����S�c�5.�����Փ��a��F���Ȭ΀R�����<ն��
�1BXHCH!
�9_�s ���sJJ}�O���JD��]���h2�9<s�J x����#2*�YD�2r�W塡t�VS�bba��DN�tsJ���ص���R�Ŀ���C�2�r�P`�I����AeE3��`�M��S��ԧ*�����z�D ��MJ�|�E<I"�i0A++r�I>nb�W`��;tA�L��u|���]��͡�⤝aȟv>�Ēg���S~��v�&�'���}r�n鏌�R����-��\�xRmh�����)��_����56G�L�-�7vح��C:���Lr`��K�J��5����OV��v���C�δ�f�3ej�������}b��3A����`ѩwŐ���R���T�S�6��MzԪ��Bb�va���%_�h����8B����ʤ�%v��)jhZ�������bb�zU<����P��0�]֎i��ee��+�y�c�un(ĸop�6�����:|�fw�'M�@}Vhܡ�Ս��a5�vW����M�%�{�=�%�������k��c�����|�W�p�����<U�����!ccf@�=i�Ӓ-!�;�?)z���[��V�?�G^����3���^�e�U��ۀ�B�0���U4j��j��^�0�5E�_�z���G�{����Ժ#K�tj� ���֑�.��c*qP���9��È���=+�:9�D �ȴ9_�ȴ�j(�����nMvhY�FN�V�6�/��sy��~3O_-�_�ڛqΘ]Z
AL�pwv��s���+�`�C �r��G�^��׍	�l��('կ�\6s��F�vj'��,�4�jT0��$\���b'�묖ҷ��?���m@/z}I�Fi4E�,G��V�.0$��C����ϛ0u�����6r�n�6Os��/U��"~x�ă��������Vp���MI���,\��Y&��:�&��C=�K����^ӧ�����@��+�4q�&����t����\ \��+Z�У�w��*�.��g����>�5m�N��k!b�o��:aM��lc��$@*����y��C��3��$���㜍���Vٞ��m���W�z�p���K�LV��s�{��'�&V�=� 6J���Jh��g(��/Y�"���	���N.��%Ѹ�
���m�`J��-\�<�`t�i���m�'�����'/�Yg���MȾʆ�פ�l�����Ax����b�X$|ʩ����d~0�Q��H]��j�i� af�"��ѹ�n�h���ݬ�M�A�w�&�C6.�4].ГX�5�ĥ�z�$�S�)��6�0�+A��O�Ϊz�c�j¥�Ϧ)�z�3���
�4�`t�r��7���SH��0����zD��V�2�����=��˥���]�R`ͱ�O���[�%�-5�E�{}%�Rð0����V`uB�z_nO��\��۷�Ć��>�"7[��;ۯ�K�{@\s���}w��7��w�y�k��O��/+b�s�W6���':����cx'z�)>�}�jpֳ-�%�Y^�`0�Q��<�@ �iZF��'sD��O�������L�B{���\��Ç�ԓ���~��7��SS����*���CK�w�]1�X�s��͕��L���Cױ�.\��LP���Þ���Ui���R�����M��ğS�ֵN�g�oکK��̘��ж��AڊW�{\����K��B���b��


�^U��?��wWޑN,�.�[`>.EY�Ӌ�$���'��C�S6M ���ͧ���#�@_�D���wS�$'m
[�F?q@W�39�Zr�뛝��o_��U��WL��V��^-O3���,-��ګﶗY^>Ї��;���,�u��%ꍤp�����z��yz�'�8�h����â��_k��ը$!�s�O���S7ט��966��f{�����/�x-�wq'������(nܣ#Z���M�E�5�GВ)QS����ᮙ�����h/y0p�Q�IȺz�t��b'���r_���Z��_X��3���}]�QÿӴF��c�;��ޱ'.�#�tu��P����̰�ML|,�b�c��5����p�{i�x����rH)R w�mz���q(�	�ső��������P������-�:=qZ=�[���T�>5�8�-�)y_�BA����8��`#���7�(<�x�V��4�|V7��؝<Y���M	D����Rt�ZZ���n��4xȠ�	���b�H��_f�E��k��L��.s�3�tl���?.�u���a�z�|H���$ 6m`/������u43_5t=
݋���4���O�r��&���`��s1ȰDጧ���~� ^�h�3�u����mΤ�g��y�4R��K�154-�уc���y�n�p���J��Ŏ� b(�{��l������9�#�}9���L��Zf#����D#R���`����p��r�Zf6~uh��7�/���&E���`��.@hy��}/��K��竂����ٴ��.��74�I��7N8�O<N��[|���>��'�y��W��[L�D��ۭ����l�]$� �9@HbD}�2|
��)S���Nܟ��<o�y��cʰ�X�~��W�l�w���n���+4;�k��܀�=d�V���,kA���-���N܏x@zl�6��B�˫��
�ߊK���������g��i�I=���зG�q��n���K���P�575��D]Y"�A+���,�)R�lj�����Z|�,M�N�|����]�魀���N�$ǌ0�7p#n,9�i�Ue�;t¨�3�ܐ*�Gp��q��HF��Wf�J�H�U׳��#�RmF~��4F3c�?B�iq#�[�p��hϔ�{%4�+<���C���Ӏ�婶� 63m��3���G���I.
o��q
$tu��^�ڳV4)�:9�J�M�z�\�d�f�I�˿�be�oi)2=Z�LqM�Z>$�d_/x�'��s#���	�� WKe�������p��feQB�� |��͛ae���&$@���q�>|��U�@~��h���pY��ѿx�A�č�n�]�4��Z��g2튶/3�'��m��y�����ڞ�H@�:W��H�8�-;X�͓jXc=�d�&	
�ΖO��[���Q��y�o�hm����Q �$̾P}g�Z�Gf21����'��G����J�4T@� �2@�_8���n'5��:��g8@9�T�-}]Q6�a�ú���9��!`���"�W%!����4%��8PrßR�r�p�(�&�T���')�+ޙ�u���Ra��7���D/1vm~��C�pF?�h�Ko�V"m����FI�QBC{_��f�B@p+�(��縗f� {��T^�[�7�R]�Ӻ�|!9P�:t���l<썥��"��'���@$K%��E�6�Ѵ_�L,��Z��b8ߏJ͏,�H��bx����������z��O�u��!��MoFC�A�<�*��-���-Q���!�!؄�^�$88����e�F�^������3;��2��"�j�#�h��n! -�6�����Ҙ<�T�&���U�_R��F�Q���I�n�7��Y: ������O�7@z���IP9�B���)�d���v�g��#�ݢ�2����3��g��a�?$KQ���+E&��Hv-��H6���2v�Z\a�����ˍ��ɝU�c}Y����G��%��BuW7��a�����#�B�ӟw���F	�x����i��x�46�Ok�:1[b�\|?���_�)e�2vy�C���v�_��.��~B&��J:�^���o�k�0H�3��Df1\���O���&֢r���s�v5����M�D(E�?���:��o�+B�`G��e��Uw+��R �����v��'�{�Lq�*�qm;ZS2�z�v�G��ޱ|I��i�k��h�/��"_�3�/��.�Ś0�W���h�T���r|��Q���;���D�����{6Jw�-4���S����¡��a�@g�SIؙMx�	����4� �^��Ӧ?EFl���4����V����s8_�SƑ:���7	!hty��]� �z$s2�>{��i��iK݇����'
=����~` Ȁ��;VIL F���V�-��ȿ���P������ˇ��W*s���X���A�>��p�R&׼��,��x���On�d��XPl���͵=꠺�;tKշ�fꞀgh̠Vh-�WЉ'���A�R!*��$���" q#�Ku9��Sb�2�Kc�0�h'�D�j��MG���h�0�
�pI��M@֝k�z��0�3Ҙ��<O��x:�����F�}bk�2;�%����a[��B�=���]`��r}�H�9�׭:s��Au�
�+j��wY��$�-�ftZWȳ�l�l�z"���A\�{m
}��C�&|w�Pv�V+t{\� �v�{x'</��I�bh�'��ۮ�q�����ա�D��w�m��J�8���L� ��ee�R���h�ݽ�Q;�M�0哺T4|�N���c��+�U4�b�,"�ZYJg�n���V��H��Nz�,��$�cx�W��zl���u��*4�c�����v^��� d.9�D���QqOχH�N��N��+rQ���n�����C�����\p�(��G� a������۞�3+h�$�ޱD�?�9���.#�5�����۞fKV,�����o[�U;wI��.���03�4���EE}pYѦ��ވ�Ҡ=������y{�6F9����D��3`��ZK��s���Nh!���k�Mȯ\�#ψ~��̊�:<�* ��e�_�_�@2Q��*%��lΑoS,�4��(55��_�e���P�=R�ϓ�0V�/�A�G�0aM�V]�}���vv�_Ǆ��X]�!�a;|�P�v+f ��*Se#��0��W(�ԟoTi&{<J�����%��2�m����_,Z�{�)��Q]��H�qA����#�4���C�<����`����3�P9��Sf��-2l��U1t��2Oխ��ئ����>�	\���i�1l,�-�G2� z:���K�b�(�g/�ͽ]e�k�V�o����߇�X�5[D*Ĕ�r3l^���ajሗ.2�}��k������*����}�a��]����DG�>A~�i �=��G�l;�s��,݌�\��	��{�d���{�6a��߁g��f�����:���@��6S\2�"c�QU��\�K�Cz����� Z�q\/��}P�R�{#�{�N�}b��\�;pxMN%�Z]U�;�MՔ=Mǵ�T�~�W*���4R�h�@��4Tp��eWC|�Z����̧.	Ե>I
�ys��9(�\��>$S���[t��l�}N�t�lD��1�p�⾖{�i'#b��D!��w��u�ڑ�ܢz����J�Of]i���'�5��.�7��t�1)$$�/���9\b,�Ю�<��R�ͷ�x���32�Ӥ�ě̈s�����3��/P!���Pڽ,,`j�Y����E�Y����ס��r}���3{�C�mz{� �����FQq�&�Bv�Lޚ^�v&jz�;bί��f��s�9�j|���9��j��-�k8��+ڟ'F3����Z�;��O��@�Y�l�8I:�4�`�-}h����(���s����M5�֓�;��UJ�Y�h��_��=�Ϋ��&��z�rɐ�ce�u�I�YO�3��o�p�����&}�&L%ת�ҥm��cL�,nF�� ��rJ�шG�e?}r��@����NL�P�V��}ݓ��U�%z�?�09�e`�]� ���ȿ���t����('k�c=��K�����9^j���O�'�L��v>�}\ڌn����h�y��ٿ$|�gCo�WW���3&�J<}w���߄]1���U>�����TTCe���Qf��C_��^�5�в��L���e��XD���#��c+����$��З���=�����m>d��~"���\lzQ���`����SC��ܕ0��-)��G^ooW�SN�}|�����Aq$�.4��o�'�������T��vy]�p4[n�����.�us��D�E_�C�G�<X���iV��<��C�U.!�@ٰ�7sj�w���)wؽ92�mPr��v��#�p>.Ƞ�snæ<h<�_}�kʂ$W˿��2�!h~����IR>�}�2�$���drа����6xs��Kx�믁�;˟a����2=���%���.N(Z7�7K^��I��RV��A��8XF�����;�:�$9*�宷�x�iqtG����뮛�)��*)��{u�e�9!���!���45�ﾎo��H���bN$n����4�Y���q0�v���A�Z��ס��&J֤�[.��x���V�ߠ�gȮ=ݭ���m@���{H��,+8VX뒞������2I\=dZ�C�.-��giY�<x�W�T{���9�3�*Z��܎om�ѧh]��:�"��;��l�ə��\^��؏}{O!�p����*�y��VQđ�L�����s��t�m�̎s��1q�>GM�+y����F����_847�آN�HR�%���F����D%B�Kd;��2�����`خ���fbe�JY@�q�toL�|��	��j�����p�J�G����o�#d�u���Q���^3Z�@��Ϝ��U\��ncgș�!=p'�@��˂�=1�D� �qK�\���)�@g+͞���;�I�*p���X	?��#Q���f�m2(r��4�|�'�DT�y/����AIթ,��xX�f�`�0��� As�jd0p�H[�cPިe@����Ĥ.���5Ѐ�y
�X`�n�w��*��w8Q��v�^�F�M@���]��R��
���;;]i�E1]��K�n�ȇ���sX�^>oS��5+�]��ӝ�s�
�w4�x�6G��l6楦`�|�[	��V��s3��C�Wj��A��^�=ً���[P@6��Z�1si���ېk_��Am�����65M��6��	�J}ͺĊ���>_|�sL���o{�5��a��,N+�+�^�t��.dj��-���%�C���d�9����Q�F��?�,��/��-�+ۻ�{G{i�"F�J� =��"��і�<����0|A���r���7m��;\>5��l9
]z��&g��7?I��$����JK�s�����.�����it=��F��޽w��{�M.��� �̏;��$ͼ҂O0W�����pE-��2"m�����l \�ں��JW�3�l���هga�8�aE.~������XQ�#�V�Y�v��.,�6^�֕d��)�b�<u>H�,}۝�xf�TY��+��T{7�.��2Y�mw��oy� u>��tjyѫ������tM��#��&���wK0u5�d�D��<_��T2��l�}b���6��]�b���3wl�?��&���m����Q�Ha<��5zHrrv28亡�:|)�
$��:)2ć��t�ŅY	U��G$`�R��c��k�?S黆�RlW��g=��W��fӓ��dҾJ3�Ȝ��͇����L�ȓ��T󋈣��YR���Ǭ�K��F�C%dOS��a�e>QH�8.�|*�uN;*~hD��K��y�+����t�v�^��U{�l}{l���f%�MŅ�*{���c���U�ߊLn�Nz��)���y��#�1����:Ol�nI�Lm��3�G�"
,�i����=\�S�x{u��cJ�b('�q�Y��ug���V&6��1��y�!~�t�o��2����'��z4ݘa�+����\���	��J�vu�1��Nyɨ�xl�If�\�ע��KS�
D"�j;��c��}o�"��C˙�����/{�x���~f�'Mu����L�N�$X��iU"�k6q�in�����d��B�dt������PZp8qߐ�`�+�1R��L��RD��qj����&<����}������nh`eկ!��u�z�
daeW��	-�������(>{":*�ֺ�ʦx������,^	6���~ɴ�'}��	�����I�r�;��p%d#V����/<k�8�W�]Ȑɇ���Ϧe�Ad0%�f�Y ��D������c�*���w:�J�ߤ�*k��{Y-]X0H[�k������x��{�J-
��m�O5^,�:b�M�N�W�����Xi�Y��\����w�K�1� ���ɘ�~RǞ�г�C�\S#��uhE��7�d��F�γ-�b�zHD��[��&,��	�&k9|���N�:��n�cռ?�[�;�  �G��u G՚F>�V'�53�,^`9uR�-�\k@G]�3��Vvamhv�j�w?w�c�av!]B����0��ǚp��O0m������=�4���6���}�|����.�+�tl���z_<uР"�JL�/%���O�]������������xJʱ�����/�A!`�I~�c��0�� )��?��g:��AUV�)b���](���JtK��|xF�iu���|��i�+K�{�K��z�v>|9&(�y�Mw��F3�r椷S�6�fӃ^
=���]��AH�=�]�w��^������ٙ�#?�;��R�ΛWs�-��Z��X��.�e��4	Z���KX5ׁ\f�0�P�'��o�wp.�+��)��p�H�OqZ�ܞ^��o��S����7���})[)�� 띦�՜��u�:��.W�5�㢾���C���Xn?s	J�������d�fއN�Oz�́ۉƈ�6:α�V���c��t�8A|�&:;��^(�䛩8{-˱�X�x|i}�qs.���`~�t	/P�C�ޠ�*kll�&�K���IrY��_��V�*����,�gC*?;|;��$��\[9��g����%w�-3rf��RS�����\����nwWh `�����<jqјzg�;���Z<��3�Bu0�C�=9�.F�#�4����p���۸
�Szj�O���giD���AJ��z���q.;������
��:Vg��T,1�S���e<3c�97W����5�y_w��S¨F�G��c��bC�۱y|un�O�3�/gؘ!���8�A:E����崴�-9�p��-�C��"��;�ɧ�+r�b�O���&ú�E	,�o�	u �z�S�E �'~�n���u0g'���e��Dا�Q��w��a�)7��� rX~&�Ь�?�;�����4�x6���>�It��^�h8�z�RK�y��]�r �vF9�.�%}F1�IL�L���ћ|�_(��\E+v%� V�/���EF{�^AЮ�+wcm�|�~���5����3�V�sl���q�pcJ�).�b��Z�sK$�D�9=� ����U܊�N!K�D��?�������^B/ul+k�o�t�>����c�Y��͒fӗ����������k>�����˱��6�rR�ih�T<���+���T�o�Y;?�tF0XC:��xPC��R���gjs2��e�6�ɒۺ^o|��<��ڻ6ј��L:6����!��X�x~���5L�Ce��V*�m�'����1�nl��;�T"�����LZ�V�H��GQ��<�Ψ�����!��@#4&�r���y	������{'b'�f4rJkн@!�l�Iv  �+v�u�c������2.Jo���iD��k�9Bf�"�CR?rCՁ���n	;�E�Oy�үcz���w���!��z�։!��7�A3F�������y��K��x��l��;�ʐ���"��;��;��r�����~��Ր��f���d|���K[&�Уry�!����^���H�t��2K=I�=���G2wD�e��gg�e�;�G�-]���q��?1��X�����=��%��,9b^Y���9XE2kS?���#��������xI!����	�z��e=��TN�O�*��i@��)��U��c�a�����.&X��%6���æH�[7��V�dn.��U �8	�f	|=���Ϲ��ƪ��gGK���o5�ͫ�}����l�=�U�G�})���f3��k����p����OϾ��L)ra����묁�� ���� b*Ӿ��e�[M>�3�!�aGҤ�JH�#��چ��}�V�ڠ6���#M4��\xAXi�y�����V�*ȭ򘡬���� ʚz��XD��y����S��Vs�4�j��� h�~� w��Ք+c��b��2�����+�_eW,�ښ�g���B<k�^a��?;���3D�k*S���}.G>M��$D�����p�F$`~?;3 `��Y@�7\�[U��^���h�+<�����?��jR(ͦ�x�����	U�Ϙ�\���KM-$�^�o�Z	s	=7�bj/�;��>�k�͕�G�l*�U�r�#0�8�q1T8W���﫩3�xݞq�6��o~`��R%�t�3ᖄ�q�Q8�:����		�,�Z�L�&�����5��?�O��Á���=���WR,�p���be��tX���j g��K�\�U,�#,�f��s��Ba�%���vM�n��ڔTL�I��l*����!9�����P��и}-��8�~��
#��̺�#������sT��ʕM��%��8��NI7�D�����5"��v�coӘ4Xp��7Ph���5/�� �ć���2D(wW�2v[�KX��'�R�x|nm����7JF��)����s����|�y����>F�v��)���uc�klx���z!�Dl7��%-�Uͬe����v��yl��_��b�!TJ|T��.�E��M!b�S���rWO��+7�[�X�~&u�-n���q��6=�4h�<����Z�J��#2�'�	/m���B���oI�Ղ��G�b�����P�I6-�<L�}�*�)�f�@��ɝq`��ƀ��pb��i�աnV�7�f�,�$[��^��j�~@���^�0�#UYqB%X]M�����<ƨt!9�_q���'qrY$�����h���6��<Z�Z~!��e�!�� U���� ��Z��q_�5�{�Z�Hp�3�Y򀩒E�٨o�VGP���8P���[�J[>Mό�hy>i!tcsq��e û�o�iI���IG�n��R����C�U�p��&�*��襤�5^1v*���~vVy@$���/�4
9cT�uP��E��`�Zn%wQZ�B�X�N���ݘn�yX�|�������!�G�~�Ϥ�J�v����ٖ���ia�����E�%<�s�����~��3O�ҙ�v�V;����@�c���+�*�;M�nQV�	W ��5</�C�{�+��sI��V�s������C�S��j�>����T�w�v��f�L[OM���l�lt�*7˧��|���B=�p��}K�{�@�\Q��3��K^vr��|�p�[B".�����*��iU�شp,����%}�&g�N�9�U$����ݿ��z�+*(ڽ?L	G�<� 8��k�6��Su��I'���v��nO��{��YTԚ~D8��~�v�J��˾�������<��[S��iP �r�Q(����I�n!�:1C����V3�`ھ���R���F$����BMണ-����ĩ�;7#�χ�W]�JfM;���يf9��K��/a5�@��6��0	dLE�)M�O���囘Ҡ;�%���d�L�}ir5@�*ܦ^|�78wV���>�>�T����}���g=8Y?���B� �h����v>؆��9���
t���������V�3a![��1f������X�6..�A��J?��D�D�fP�Lw�价������{�u��%���dX�	�[�����Ý)�د-��e�{�ꄄ��b3I(�c7����+��n������a��-O��V���З���+���a���"	�L�@Oo��m!�]�o�^��n�V������E�rZ�UN�F��#N������ύ���CRa���)#]�����˙���=b�����۱��T��Mk���{萺:6�"B=�\��z��@�-1)I��%��|�����z��k��ge��q��qҵ�Gb�{KwW�y���6�qxz�I�I_���k:�tv��N�8U ��N�QլJ>y�z������e���pm|3�ZM��0�S���G�%8�����~a��G�Kv��):TS4<�	p�v�t�1�,�_�-���||�Oq�h{�ϛ�oԯm/�1K5�C6��)��!�Xh@�nT�?�=��_>��i�br��V �_��Yu�A�F�lOSs~��J]�|�ⓁdIm���"[ev�ߞm9�<��gO�S2U��5���KG�7 +	1%�R(���B]��~�-��S�<��G����t
�+$
��b�c\����ռR���AK�̈́n*�󮱵K�H|�Q�Y�s졹�.?�n� �R9��*�Oe9�N_��oB��?����B�Gf��x�'��w�~e$.��Ưlb��7��	^B��
J!�g��.L\xA�2ojatA��%��ʌ�\����i�I��������a`L�yNVtȘj�h��74Lc�O\ nA h�K��x�J��Ç� �D9��V�l'���Q�:�z{�U&�?3:q��W�?,0fA���M�����2�WQ@ֵmtgL6�`Cᮔ�(��� N�H��:�e�4T4�>n����>��F����[�P�A"��N���|�'���2�����wH���ϟ;1����Ӯ�ۛ���Y�g3y������I�� � Q=�[�gHstk��\93V�^s��T$���n�ɘ����
����%($T�#�(FW��F��r����T�-a8]Rs�ӻR:l{kވT�U�l�I�8k�M~ʞ* �~�dn�]��m�O�w�h����gtV��
l�ig]ñ&|��IK,���dM� ��}F����@�UP*ؔ������Sjj���rN���N�d�T��pW�O����*�5��c�â����QDP@JAR	�F��Α����D���ib�!��$��;��<�������>g����^{o�K�/ ��p�n�&#��;�V]w�����n�T�n��S��7�M�J�H5������նGo.1Z���?�C����~9_�:�TM-�d�H��$�m}�[J��
�z�Id�L��h��ni\s��d露 �m�.&��8Q�>��7����h�ꃜmY���C�����ӏ{xU��)Ȳ�I{E�󉽺��L�� QL�XwWn���F-�\�o�4K����2c��Z�5�i�,�T�kڳXJ1��F�C�[�&��C����֛��+�
�	��y}%�<t����k�R\\�^&b�0�v9�p��^� _��̒��KXf�[��a�.w�5k܎%O+y//�l�;�m�޵�"�U���W�FtJ)\��3��I��R �,	f���i��mޏ5��z)���t�Ҿ�����"&l�z�:5�\�(*�`�W�F����T?�SQx��Ӿyg@T��t�<.�l�dw�6I�+��:J'�۫�S�V�#����t����Ώ\�݁�o���&m�h����ó큣o��ioI^8"ޠ�q���#erfhRV�[K7u�v�H	�&��7a��j���lMJ~������y��̾�o=%A��q�]�^%�*�> �65=wy����SX|�f��=M/Î�-՜�@Hǟ�S�����ѣh���+�~&�g��~a����L�l'�����Z�L;�I�M54w���f���W�u<�Ϧ�t���pG�DW��o\x?�B�bO|��^J$����t}��4D���d�~�[�D�O����M�+��ۺr U��T���B-3���؎퇣g����۸�j����,`~��*�a�C�W����}���M�C �e��E��Tu��q~���W��v�A�I/̫P4���x���u�[o��K'��d�mC�����[X�NKb��V�_]�r��F��Q���1��cY�����Z4��8�/'��8�0����-Ѫ=DgMX��s������Pw��)@��"�Ï�؆�O��Ɔ*U958'[��o1�7*s�rbп�/��ر����Ľ#⟬8ԍ"ӝ:�_�����h$�u���ER������Z��^:'��}Ӟ��~�������[�7MI������y��n�����e��;r��F[����D+9ܓZ�FW+�b���^V�ֱ���|�8���>�z�k.�:΢�b��2�0i�;���H.�'�
-'v�N�j��Ή!�W��dw�����1�w|��-�����D%r�o���dp��_�'9�'�����"�M',8~iZ�,N�FQ-��w ��h�� �0X+�
ƥc���)�^$��N��l2���߸�������Jg�H-�9��#��i���~_�F����f������e	Q��v�ʭ�mh�r�5�3���EC���{�a�gktk��=�-�����L݂�`	�[5m���t�'e1�����l�F�*b������dJ���a�=-��M�Z}��2r輰��|�nw�Y�py���&>}��x�m��%����Al�B��z�O���t�L�B����i�nOm�Ƴx)��o@<BZ�3l�g�K�����W�򎄋O���G���� Q��5�਱C^����X?@���΅&�	�j�-"��C�m���t�FI�
�ĪK�͵�$ej������F����)��<U&��^�%SL�$��\�=���^֠�D�-�]�Xţ"-m���3��S�bه���G�8Ḽ�S�r����lި?;:b��7�.ǔz���3ti۔��?��=P7�}&n"�{fjPk�ݢ�\�E�v-i{�r�G�I��	���W��-�c�Ddp���^{�R�&]u���ˎ�K�!#<��Hɑ�-Ȓ�Ї�WuI�5��~z�f)ξ���� ȵ��n��I�/�/�K%'�ҕ%R�O-���a�+o���ŋ�h�ܱ��o~!���R�r(����h�y�S�{��b�P��+	f��Dv o��c��OW�qv�Ep\��[g�j���+�EF>���}��*��n�5�ۧwg���rw�>C:�VG�w']�F�ւ8Լ���� ��y張%���cn�2��F���@NA[�w"N5f҄_ԶT��,Mz{G2�-[���9�m^_l7z�{��.Q����g�+��̭��y�nL��Vх3��֧�9@���d0Mi�w��3��$گ�LH�d+Kˁ4L�g_J�}�4�˭pM�
����e緧�dBX\hr���u��"� ��Px�[j����6�R�7K@�2z��ܐ�l���Aa߳WEפyM��||����s��y��,�`.���H`�a;���&?R͸tOa�!,���6,�6�8�L�{�;�K�����o����U��c��$SY��}O���˩`�AR�{�������q15��W�H�J�Y�)j8Ơif	�ʅ�	�b>x�Y�P}T��֠CrG�Ϛu��~����qLx�,���
��}����v�j`�`Ũ[��G��qQ�ب`z��uӄ8����{e�@�K��]�.���M�����mvw�T8��SDJ=�I���xϷ�o�;����}�.4�|d�R�|�#L�:ܞ�(r�[�� �V$���g[���� �d�̽�W��d7@���4N~�|��&Цg6�A2PC6��� �q=#���E��� ����8��7��,Iz�>����q��X�t����/�T�1����I��Zf1�s�/�~����d�:���4���a�h�Sy�����Iyw�Mx}�U)Mf��Y�ԥ�?쭣�N�˕N#��v�/<Zo
����LoDtQ�p���X�QC|���ŷ�H�rJM~��#�;ـ}H�fJ��M�6����:&7þ���&���!(�n���������U��CR����h�O(-�r`���o��c�V�����D�өF��%�D�ʈl���n�s
cA	��6��8��:8�F�ܯ0�߱�q��!!�'-�wah�c��J��j��VV5�D᳐s���K��#A���=E��7��̻�7���-�$-��<;��w">�t�s'�	�q9����|��ӭ!�-���\c�']U��eG�pPs��\72�����N�P��I�v�����m$��k�|�_��G�T���TD*��*ؽ�0��T�JY_Zx�����:���j�L7��(�scaQ��k9Osvq!'����;<����.�m��fa
K�����)���C1B-���	ub|�p)X�hC��9Ŀ�r�8��`�j/g�����ظ\���s�Ol4������E����
��=��2��E8�Y:�cU8�&(�LK<�9���n7n�uç��X6�� �/�z����I=�`D�?/�]R�AOH+�օ!JyCe~�@���U�/0�Jd8p�Kg<<���Ϗݷ��ĽV"�>��J����&�L��Aiâ�gK���Oy{-I�	�w**��%i8��r_��Ⱦ8���K������tk)JGz�%:��۬C^�2��(h�U��kLh,��eY���ي0� �~��8\�dW�/Z��%���^s���~=,��(G����VUJ#{.�n�#;HZ���,�mt�	Δ�}q�I����3�@@�������}���Z�E wk^���2�H{��]W�6��iy�O�9��p���oZ)��-��ǵfP?�<n�տ]�$s#�Ȯ��q0�(�u�'�|����щz	x�j�)��x�x��S�?vj ������{d�Q��Sd�c6��x@_��Mg�	E�TZ%�~EeO��/d ���s�l@6fLa��������P̹G`�5����+l�B��0�/�B�߫1�VC\�ȸJe5|���)��faҲ�9a�S��\�*��F�JUW�e����9N�����$x�ӌ���%U��c��
��0�Y�����y&#���X�=['Bt��H'�-jf��4zI���f[�W[)���������U~�Y5�Fn�����#w)��C�B�Q���A3�h�|?8�%������ݽaӐ�K�?t�&Z��G�&�4W<����g�}a���@u� B�]EcjLC�C����H�D�R�+n��{�\���:E��9�m嬥&��!�Z��<�[u�{����$��}�Z�
�P��a�K�%��Z^�*��\V��/,`������z{ �����=����n�j����=�)�%�M��Vur�z1Kәrq��Y�OxĵR�!|7�'�� ց7�".~��T���-�$�;{�ȣ:d�`5z��h��MP��_�g��"$�U�X�S/�n�=^��j��j%�/��o�c�v�뼸4Nƒ)+=�E�A=��ba��|H��BM�Z�e�53d��S>�\ż���S�^�9Sw���#7��=%�F�<Q<aoۗ0�[2d@�M�$$4v"ė���k��R P�tϟ��ꁸ$_Z7��i���^h�k�nX�����I�I]������Ȼ��ֈ�ɰ_�;Y6��n�ʻ3����	\n����������1�\�e�Jq~���jB+�D���"{��
W���J��s��/������W�qBGme�Q��7W���u�Dp������p�Zf�P�N@y��3GY��A.q��T��q�%�����BM�]��j��ϫ�,�Y�F9�~v�y��l:4�M�t�b��_�=�(%������}`�������(�����T��q��2����G/��1��Wn��L'���jz�_�b�(9��3���/hH��q+�;Qx$J��O�&,\���Q��Ҩa��>����v��̢ח�s�:D��}D�x����.B%����l�Q}C{ ��d��C9����7A���K��8�)�z|
��)��d6�ۈ4�s��r���Y��ဓ�23����
9�3� b/��ǅ�1���l(��A�7�����L�F����k��z;��/Gg�x̣��?cbW��r���,zEkz��I��px/��]�5�$zM�F%� ����s�A���2���ez}ݜX{m��K(\���?�0�'�}�f.29��.\8��U�\=c4ut�T�c�0j��x����X��U��
��=�AT�@���c���[��"ݬ��M�0T�4b���]I^�K�nS�?�0���cN���a4V\ӏkT��UŖ�oЂ��㷍����,�����S��=ψ�r�N/#9'����3Z����d5�I��
���W���[?��PXC{�:r,a�R����"�Na3yQum�{�b�\�)�B�x9�z,=7�T7�KNp�JDbb��b�x�洰�����vD�#���B�V�8�6�À��[a� I�kq����;k�gQ���ۏىhO���;��:��ɨĿ�S+��`àQ@*�ߚ�EtǗF���n����{L�AD���[a��"�o	O[�/ �o�9����	��A�f����d���+?#_t��fqn������g�Ʊ٬%9O$��*�u���[-L�*]� �d�H��"!b��3�C��먿zZ�ڮ �3�V׼Jţ11/?.jjD���B�z����=
�4+*rn(4Ϸ�d6�7�����K`+u���������F��&pw-3�;R�f��i�H���瘠[hb�@�q��G�&�:�_:�� 
�{��(XQ7=L��<&�m3È=UԙQ�DY(#��CZ?�ƛ��Q�I���]w��A��g]A&���_y���;"P���)�N:6쟫�$g�S�,*'��f"Ӎ���l���sԩy��̪)n�{k3�2�-���x6��B����Jn:
��k�55/�R��0@8���ۨH��/KT����>d��ցd� \�@?��n�o��V�'
x�Tg�5J�M�<N�QAw�\\�De���=�N'VM~�A梪C����a�c�@x.�##�w�9U@/}���j6�q������Q���o:�n����ϕ3Jh(TѰإ��U�C�W��n7�/�Iٽ��M-3B�(�?��O�R~,O+Q g�����ǺĪ�j.BH�/x��x	�(����k �����ez�Ż�q�Vl.���K������-f���̰�k�:�Đ���� @#q�/`(�РRL;q�ϳӚ���
�_\2�����ql�B�:	�:�d���y�G�U����H�C4����ʸ3�4��ޗ��7f���<�T���r�Qj0@�����6((����Z����h�3J�i�Uv�6c3;O�Q��ɒq�h�<!�ʿ�:�G�i��M�����u�W6:d�Y�D�:���"�)���TCkh Uf��)�"XpE0z�q,�lѓ�J� ��`�Jퟨۿ���L
 �1��w��eg���#nf���J~�H���5*G����i6"d�}B������
3U���K����6��,'7Ξ�F�������rO�����?!Ψ�N&���k�-�U6�<��h�O_W,�0~EŽeE^_{��C*i��A�`�Iw������z1G�>$wjQ
6����g���@�}p)y�{�5������k�A���{@���?����d��`��۾jf���{�A�V� `<��2^�r�Jλְcf {�v⿿?y�Qs�'x�}5�Zd��sv>�=+��uG����Z��p����� ���ì�	�s�{'I	�le$���/Dgss�"2*WO32�/���y�l*�lIX��a_o|<���I-SG�K9_���Te�l�](C�a�l���v�lآ,s	�~U�=_%� = � ���uӾ���Ռ��f�$Ѵ��#C-^��"�p0�*��X�Y<�LK6���v|r���ĸE���y�}���%�t� �a��l������0`P�d(���O��q�)o��t"�<�q:����A2 @Otl����ChG%�&���=����:���VI��}����|4���৭Swf���R�(�-�T&O%.�z��쏩�
B���� �~i��0�>����	� h����N�N��Q�&8+H*j �!Q� �^�� Ӝz�j ���\�5�rQ��'!��7A�'.C�{L=�.\������ ��K�Jw�aR*��ڍ�-�<�!S~깚<D���a��O�� �p�-�a]���g�L+�G�wq9�%���߲!z���ZX��sjX0x�A��B`$0Z���`&�R�p��e������c/̆K#���gL�m�ŇUh��\���s�ل�S/���x
h�R|�T9�9�~ݔ1k�p��D��OU�����m�A��m��e���G���w������0+�z�ߠ����O��Fr�����5w�t����\��W�D����[��@|���JU��:<{�O5��墎~Ң��~z�o-|"�@��D�z�{�@��X���u3���&1 �@���L�H]�ss������	Q�v9{Vx�f���;4qh��Xb�� 8ė��G�'QA�4Y���B\�B˱H�},*�\�?�b�v�� �ӻ���c��w�6��4���H�s7����_���s����� �x�0�Q?5t�#;����X�,p��q9/w ��$�Yp���:���7�M>?᧏�������&�mq��h���K�Lm�/;?O���-;��,��c֯R��[W�)�� �+��4 �䀦D�B�9;b���)�w���oQ�ZP_��� b-9���p:����r�Q��\z3�N����r��t9n�q�����q�@/-��J8��9��U�^G���5}tGt��i� �ϳ��&��������;k^ir�$;G�ql�^������Ա��϶��(�h�f�!'6H��� �0�o�%��/G2���r��쥓@|�8:�KVSS�Xdt8;6�.���f�M���f����#��^��{�a�������.��X�?�cz���CyrpT��>�{�K9: ���kArQz�����"2A,�|�;W@���7�`&�)�>^����9.H��d���v\l[]^V��i��@� &
-yӿS�-hי����R�'3B@?���m���kU��0&�X���h�BN�1O; ��B��"2�2/�l���z����H�O�z��0a�i2�7_3d��Ц�B�w�2�2��Zeӄ������C	E�
��^����~s�'�l"�t����F�m����$ZQ�����"�r�F�k.=��<y���Ta�|g�^�ċ��銶��q�W8�=�P ���Dk7�Ϝf��z��V���)���i�]7�O�s[�]�r X|@����D�o�	`ܤ��8�ߥ ���������n����sv@ԧ'��j	����皵��d�����{�:M��|/%�6�O�M�b������7�m���܉�%_ڟ�6��-A<u�^�v-f���Н)̲[��~�P�������#���Ωaӄn(�ڽ��%cO(��b�����w�s\�0��9)�i����[�=������	��!읃:#Rn��ƽT���$�h��K���VbJnx��4�n�9��[]x��I 翽08ts�}e��O{)�%L�#W���o�R�o�D᫏O��HG��;/�8>�J�e�1��[�h
fҤ�:��Q�6m�����y��J���N���}��2r�#�ź;)B�/�£�����U,��͏Ҭ���A�����}��Rx��P;���٬i_���.7>���qM�z�0�ۣ��6�؝�x��(�|'n�\p��+�
��| ��S�Jm����Em֎�dg�g�E*���i�v��S�tM������������TQ%`ذ^/�--�^-�0j�qSD��Ɛ��]���F�/���K{yy�p#Xg�'s�U!S�`���	����qs�W���|�c9gꕡ<pf��ڱ�<{-��|�s1�9V<u/��{��݃K�TE��e:1Ҭ3�����É�����ł�o6D�����Π�����rb�͇�-����#`�>Y*�:�����v���{����Qk:81.�G�)dI��&�������U=��!H����J*�,Ü�Z�d��U�]tGn�`�qu�K�~:^3(�iK��hy%�?Z�%�����t��8Ё��/�(���Q�*6�,�u��1�m}-r�C1��y�|�X�\��k��HK���ޭe�{��.E��B��䗛�J�5���I�`M��
�z���j��YCi������>#��
1�u�H�@k�TWjfc!d ^���2�6���]���",��#0/4��KR�	~���fӽ���dcj��%�J>$����(oz�R���$}�U ;_�r�ޛ*t#^�<�ՂLik��3���S&�E�%�:��X̼��w>ꜰ��>A��B�恛t�3�~ᠹ�I�g�`,N�	+1�B��;�i�T�C��6/9*M�`�b�OL��� �z/o�?!�)�:�q�EY��Ch���\���4���F�@*9<�x9��@�����n���ݞ��ڳ�Q�"��.�j}�- �&�>�����cPg��s2��nH���M3�~l<�������\�::�"#�*��IH��������q�WᲑl���~���"��e��ly��+�$��g�nOҖܐ��~=�q�	Mѭ¾*۳�%�\lӭ>(��-��ĸf^]*���wŦA�u�lb�1�$�U�M�"ϻB
�LHDӷ����KQ��:�8�~��R�/E���m���r��.3<�Z�w�o��~7�(��v�C�5L�=	�^i�G�HdK��,s���������w���A�"��O_`���՜ ��n��j׸���&o�>��0�%t���vUS�s1���ɆM��Ns�[Oas�Jd�8�������l;'v
e�������6�<x����α��rO|�Ǿ�}	��W/oMߪ�qB�
���)l�SE8S0@�*k�����!4��ߚ��/�
bk�>���/	�����
S~Bq+QΏ�kE,�~���x�b�f�M|!���e並}�g����uS�Fop�N��T{oT����-`A��(�"lvFnT�0�؟�w�}}K��
���h�]�̽�׎1W/;<E��Vⵖ�t۹E؄�����)�E�&f�Pg�����[��zN�~1�q�b.��"j������?SX%f7����.���N��m�W({�^ܕYgCkP/B(?�J#�3<uB���&��E�ر���̔��,�nՙ�z~��K~F[����;�Ćy@���������� �K�hBn��s��=e�{FB$���l�x������B�,�%0( d�z�I�������(��n�(�,�ƹ���[Se�V�^l�k'^|[oӵuR��8��6�1u��]���(�(�o���c5H�=E���i�k;�G�����hX(��7c�X@_���Y�($����u�#OA��[�� �����+E�n\�A�Y���{|C�'�����%���O��NLM̨��C�d>���hS��4= �X��E����gr��IU�,8�������ոK���h%	Wo�%����j��Y}5�l�ҶU��>v�7�e�.C�J#9�F���R��j�������!�8v��CW9�kW-�%� �>{�b&q��#%�I[��6�uq�e;tLj��,�����m�·N�~��=^�
4o����X�hJ��Q�6z󚝪�FxĴ�p��
,�٧��t�F{�o�.K��b�T�Z��K��l��*D9�:�K���.AdQ�w������ ��H!M�C�<Ϥ���d(��+��>�^Bn8 z�_M��n�\�t�dp��!���)��qa�8��Q�]�a]4SV{} c�9<���*�X�j�����$�tp)L믅/�����^ h
�Nɟ����C*�u�X�Ĝ���{u�
o��;��5T��[��ҏ��4V�
2j2䪑	��eF^:�~�.�?�s�x0��=��௪�Kq	�H��(;:y��h첋E؈E?E�=����Ƿτ�ƫ�.65�	����\��Ĝ�y6��6�O;M�u-��ع�K)�b��u����g��U~7Fz�[�W"��z��5��|��\���#��2�������Ї�x
��6m)�����z���Z�O���,q��g���FP��iy��%
jګ�.�My��7����b��k�/�ٗ�Z��65g��xe�t��ce޹y7�j7�p�H�^�@�TE�ի���<��@���֠:��r�V�^m7`��*j��%�_%.O ��7QU�+T]�r@�IT�A��SH�MI}7Y������LY)&�!k�,���W2Qa�U�0�ח(R�8���*M=�ч�Wȣ��NZ�<W��#�b���)]� J�����`����z3�WϠ�����]����d���x��G����*jF�6fgU$#Pd_DΛ��%��J�`��L��Dm����~�����z����b����ߜ�R��z�駋Ҥ�K����xصǼ��������ݣ�R�Fj�NWغ�r�uu^��p�=��_ٞ�7;�/�*1_�<�8<��{�0Tѩ��;Z���<�p���K�����q��r	������Ӑ^�YA�<%
���ң�I�K1�����aw�w����۝�+qPz���f�
k��i���Nj���=�)�-����(����B�{rÖ+a�p���%ቻ�&>r����U�l|��r
�y�*U����bN��T�'�bi�%Fi��Dl`����gowA~i���$��QG�͵_��r�Ʉ�2�dj��H�{��VXI�,��N�6�u-'��0����4���SXEe�X��R�m�\]sZq%����R�,?��𕙖;�[�7`R9�������h� w�L�m""}�mu��I.g��FߨhQ��rbP�����}%|a��9���H��q�c�D�U�n��M�>L����Q|���ܥ��D�vMc��#7�9�ر�Jg�ǋ�&��~����)G~�O��<�\����T���0jz���9��eӺ�s5i(H��������m�;��7Y��d���إP�8S�;9e�7O�{>�d2T�SP���{Y��>��~��c�{C3aoN��x?J�Q}�pJ#a0Y��Ļq�h���������+�3�`����T��9�݂z�{s��=��ݕ���ν:����~�S�,�Sg_�6��W��.���o�&ANL��Og�WË��YIoOlPT;ΝN�+�N������6���,���V�Uk$;l�Kc��A`&��B)f"�;��_6�s ��/�>Y01!!fb�^���T��o���r������~�kL���t��Oh2��jM�	�	��Tv��{�|C��};��U��]i�CZ��2-Y�ЊT}̴r'�>P��K�� 7Ks�3�ۻ�z�\*&o�vn���(�H�#!��+��C�ƥ���yX-�!�_�e0#���F�2-�jEg�TR>����\B�S0,3�Y�%�.jr�4�����3�/ߍ��:��Ys��s�}�H7gi������4� �^m�;ݦ�",�ư�xd�s������[�̀Rx�� l��� ��`\�n�aK��Si��N��)�V����V<���o'��v��<�l%M��!e?���)sΎ1��4�o�Dp���"k9եlɿD�bL�� X�,1�~	��/��u�;t���(�H����7��Lw.�������y���18YhTŠyA}�9��7����)�;t�!�K�$3ˉD�;���(*ݚ_q
;��6'd��Z�l�Nˉ2Y���}�i�����Z~����K�
�8Kq;�(��E~v�=���Nx
�/ߝ�����7)xރeV@���) c���S����g���iyt�)�k���PǗ��gd%����GIK+`%d;o%WD@5���N�b���7�7��Z��w\��T���O��P��f�붰��M�d%Ak׃f�Ղ�������n�b
#ʣ������&�����#� ����9V��2��/܆Z������;�#���r��F����%��-��^{Xx�1D����:$����Bl�
Mi��N��i:p��SL��?L9���S]� �40`n8}�I��ס�bz*��Г�t�q��r(r],�_��i�*nn�],������M%̓�����4���T2B5ۋy���0��Pn��xKôzK35/|�k��	58�Y��&Ll���t=�X���ae+��ث�չ�-@v�~� ��D۩S��P�/? $�/}o������p�u��+땹��D��2�h�C��zb����c����m���nn�����3��q�IF�Bc���ʽ��2>��0ެL��WY5 ���(K&��c�`������v�m0:�i�`�7_Z��������e�t��Tqp|Z8U�Ʊ�b��=٤�δC0�TCW�NFK{wL�k���zțVq���F�%�O�s�H�/���?s*�;�a�m��;-b����7�-
�>�J [6Ј�k�#ܶ@��M���T�*����x�2Zwo�y>��S)��k ��59��u߸4�Wة��.`�u�2c���p3B8�w��j������zy���/��2��j�O�I�T�/A�E�e����f)����^ d�
M��	�1	�U�����g���]|�����	Q�����8�"���������V��p��r �ma_�ի�u)
n<�U�i��>����y�ST������-OQ�ǟ�FĀ�����o�ޱ/z���*�|���,��R~=�*]%)���7��`ms;���]�hUخt]Z�p��~
ݪ��L>�S$7J ��m�.��ꧩ�?��_~}��3��Gm�LT�*�����9�m j2��3�]{�ZNɭ������p9oD���x"M�C�*�1��\��N���������Ti�R��p����')+!�O5n���#�h����:��q�!W\�0Fj��M�>(ox8�m1�>C�!|�ޕ��$i���b��k����5�jH��$S�C���\��C° �%�) ��5��S�4�R�\�IF�W3Er_	�{<������Wai�����D�q�X?��s]8g��vr��a˗jT�up���S{		+O��J��Om�6���������/;^�Yg�o�2����&�z����%���(�P[�i�4T�N�t"��5"��P��k#���յu�א��}YW�R�.Ԛk�]��V��3?6lS��ymN$�:��S���S32�)1f��ĖY�Le�|�"����$��
*���n�����Ig�3���[��L���s�(�#��1��R|Dҋ�KM�8�&��hKـ/j�P�n-;���P����@ˉOo��x��;��s���u���D���iK�|�_Z&>�n��!"U�/!Zp�̡^R������n��EGB诳~#�t�ۼ�ڞ���3
��)Ӟ'��f��y�u(�J�s�7�b�W�|uʾMx!��spl��+�ow ����D䖯�$"�@(�]�Ԫ�y�����)+��V����k��G��V��[�>�O�x~�7l�f �x���6d��ַ��Oqͦ� B�M9�A�&�F�U��V@���Smw@��uF�$�[�QE�m����d����S��3M�C@����A$�YW{-c����R�4�S������b��>EB���9g�%�;�"b ��m>^K'��B{9Sތ�r,�����d�0?)��Q�������XIp�B|} ��ޝ��t�D�bC�O.�~B6Hb8��C�&=��F^Nt.���Ꮗ�L�˻�\�=�S��ʫ_�c�����v�J���0 ��u8���s� J���;V���
�+Hx��'�/���u����a[�dr�
q8�#�$�f�C���#MB
~��:;�'�&�����A�i��pջ����C=�=���;�.A������9�z��r$u-W��Ia[2�h���x�-.�V/WYX�H!���A�@x��Q�HE"вQ0pe�~�J��-Qk Yg_�ۣ�'z��')�Dd�E�k��4�X!����o�)�����:���5��mG�H��
{1�]
�d$����{�9��Z���X����D Xm�T{2��y��$�F�䛦�JL�t�q!�r�l��!��y߯�&y,;�I���K{#��S"ױ�S񈭻10��Fw7�\�q�P3ul+k�>g����a��ѓ*j'[rmlw�.`ت�G�1�%l��6�w�#�a�Gh,G�������[)@?+~%�����c"˷�ֈ�,�j��
�7�f��s5ﬖj?�����Y	-���k;��-`0<�K�>b���N6tP�foE�ܡ/�?-���{u@���hI��p��٣j�*�Vm��S[b�4�i�����Qe��A�7��(P'y/g X���Y'D7���R��}�Q!"��I�;�����fZ��$�	9���d���NH2�&V9�˅2���V����m#�
��;��GKߛ��1�7	�}y4��J-1���K�x���?���_=��^�3�ƭ�K�K?z��!��I�F���ѕ�4�o<�:��^��4Xщ��b�W��ӄ_f�v@j��9�G�@�����l�ߺ�	������ߴ5�Ba�e�T���f�D}��ʑ�۞g���/���y��IW�Z�&1�:􍒧2�̟ӄJ_��e�gs����{�!I�x���=��a��l)jj����C��e��o�a]c�܂�����$�����j>I+��r�^�T���'~h>7WןK�Ap�S�AA����2
���+�� `��� ��i}� 'g��6@\��8}�?Z�����W{�aj���<{-`Df^:��ߗ��GI��	�q����OwcQa�%%%�G�?pk���B}����'

t�cQ��ז^म/�I�����	�X�2}��k6`i��e���l3
^Y�u���J�0j�G}��ԣe�|�轞K�Ӓ���T�[���H�kk&A>>A���'����l��m�xd��]6���D/`$]���82�Ȃ��-�_�90Q	L�,#o�1!F�		��4�r4���jjTk �B z��G�<�m�p]]~018�K#{z0�wv��b(��>*� ��3�z���D�K^�LN�u���L��%Ɠ���6���_������w��ō�������Pw�,we�M�dX%����ꞆZw�: U��c����ߍ j�6g�V
�06W8N�Ե��EQ������{�ը�z��6�._B�l����<) ��-��VV��$w��y�<=�xEY��"/wq����?�ћ���S].L�s���E�ҳLt�m�s��]���cO����DH FG�L�/�`*t�+Ͼ6ӑNf9Qa�P��2v1�E�����������un|��,�{˫K�ʦ?�(���C�=w�Oeeè+p����D�Pp�O������%����ܢu���Q\��#�h����qP��H'�I)����F�F�,�[w�:�����s亞�?Q?G���:�˝����9fy�h��n��ν�n0�+ܓ�����ɃN����l�V�_��dؽ��'��G�U�wCTB}��e��6�9ń�I�E�J����;o�c�%l���Tm��y��!u�Ն��e4��ղ���|o�=iȓΕ���QQC��Y����I�o�c�>��a܈wݳ�N�:&|n/��a���#%����P�ۂ"k���x��:/�\��|����������Gs^�)땼��[u�)j�FM�h9Z��(���|�������!i�$�i���B�˙d�Ϩ�X�X�g����_T�9�^ڒO��!�Zt�v��Ǜ6��������ݧ�V/S�Z睔
G\�F��J��9�*ԏ�Z�i�fo�Ϝ:>���F;w�u�<��a��K���c�{���T�6!���e�������\U^�G�+T�
���S	��ieͧټ�aŧ\n���W�u��'�Ss���7��SP����ω|���̩b��������lP�t��-��S��7����gf��|6Hrf��a4�/�)V�9Z�!go�Ÿ�1nf���G��-=�0��p1^��A��к��`<O	w�O������r.�MÖ��0%���=���*��Wݵ���u�̘��Sՙ��Eg�EQTQI#3c��S�VQ���UA!�C�ִ��S�,�:$J	��S�cJ)I	�s��I��y�6ϟ�~���k�����}�}�{���v�W���z���������<Y�-(�-j"~��!����R����4�s׍Ĩ%��aH��t�|�i�7��7塜?��m���a֥��9�Iڎ���]9��������v���;Hj&����Z�.mg��W�_�!�/RXt�L��'�[��k�m��ͤ��S�����"f�ػ��ɲ���o~����3 �K��������x^�W;��->��X��ן���6���ȝ_�rӄ�-I3ȅH���=Ц[p���6§ݦ����r��q���>>g��[���a%��(���j�;��qX�Ґ.�׳ܘ��̳$ڠ�s��J�ݤ⥖&ޮ�[U�'��G�_���"t3��Z[�3GFY�[s�	��#�۵����G�L���^�Ll	�V�骴�ڞ�z�:&��O�n0e�5��y=���t�+z�{X�{#<��~F��l�c&ux-U\��k��N��.�}TgC�h��� G�[5�x���r ���D3bc��4B�.�>�0�b��4H(�?�I��-��臢:H/���$�f���&�1؍F��4|��.xt
6H�����՗�](�.�#����,�y�(N�]�c箾Nd��i��U-zB����&@���*�(K���2Vs��K�z�Fٽ����֝C!w�_��m`8��E��3�ؙ�ם,��#87�)�>+�4*N�~�@�g��-�KMe�r3gֈ3����T����Ń�?[��*ئ8�ʪz[�x���z���DK|�|��ı�;�����w��q3=�R�K٥�ՑRL��I��q;Oڔ�L��6���Z.6@�k��{PjH�Hj'��s��'^�L��s��j�>s�U��Z�/�X����j{�*�6S���@6���/
�L�&2f=͡�u�M�P�E�.a'������'0� @u����s���M>�k����L����H�.���TKnEQ14ec���r"�� ��8gd�y7��ykkw���0lΙ��7��~ct[8�&,�59m4��S[�Ȁc�n��K6�-3>�ٻ�|ҋgEԣ�I���������0 ]Ac�Y�и2�c�\n��@��^ ]׀jn�W�$ϓ���Z�5��e�1����)h%��d��$�������Xo4*��k��N���N4�U�7|�H��tȗ�}���|�p,ь�~���z��;|��]����+8��		8a`�L�EQH5�:
;�`���?+^.���<�R��~���x'�=��~a`>��Y	�i-O���lPE}Vw{eV0;�j48�f��A0�l���l�k���?O?0�؝Ѳx�|�{��\��ނ�<ؙ����?���4�q��a����V�Z
���a���N$�%��Q:��~Vl�����l_8�=<�r+���U�]P�����e�c���|Fvc���v�hb������2g]��s�`�>�S�$����W�{_KcU@��fǄ����9Ƴ�jG�I��l?� �qi�X��C��Wϱ:!���V=]��7|Do�0y�|ͳ|5��HI�X8Ӱ8�=O�G����2�a�����m���������b�Hst��vIb�Ѳ�9�C��'w�'�P1�̘�R��rm�٭�<�
'DK��	>IIYY���Gh`jC	��ղVI\����H����<~Y���4��`�w�]!�t
vس�%��N=�zS�����I���e��k��hci׷�bI
���$��z�XӞ��:5̠k��G�U.UѰ�hW���۬�q3�������n���h�{��33җ�I�W)]��?���5P���)�D3�Y�a�W��@O/3K<�������s�x��j�g����6���NL��E���2�U�\��<�k Wm�q�#�>�(:�ҍ
=Shs���l8+Y3�m�ź�+͖7��NS(`�D19O3������u��Rw&���Ly�� b{َ9/R�C/ۓ��)��e����EV�^f��� y7GP�R�3�!��"��F�1�q-S�K�ǩ�����I���0`����g�e�E��ɝ_��?-FI���ŅzkD;l�f�x��D���j�!����4��`�I��L��fRX�^ї~���[x7}���-D��]�Vr컣�	mL�[Ɓq�5�V\��j�/z��#�⸁6��O�X�RS4Kp����m�|�C�5��/W֏�����fZ��v߼f��OVG�>�"�5�i`��ͷ�`s��8P�)>���VS]�*����|�y�94��Hz��w�ݐ���	M�ݍ�w�>9P�'�22�g_Z��||�	(?4n����1�A=��M��{���b_�����cBӳ�h�N�폯g?�+%��Y��G)�D��xC/�PA�e�C���	���`C<��H[K)(��H�OٜX�S{�S��~1�FW=�IƯR�E�lg JZ�0��% �+i�koL���G�</Q�0zy��5Ѵ_�b�9jf�5ð�L�o�n~�o��c�߰��z"rs]��3,�mZ:7�������Fq�M����#J�gg8k���={-e��0�C�f�Q�[�'�$_��\>H�v{��0������\���!����S��\��*��Z�S�?@:�jm�L�0 U��ȯ�{��P�t�V-�T1ڟ���Zp�l�W�(b�&Wc�����0.g��Z���dӼñ�ѽ���ʮ�F��;�=��r�T��P��Ǚ���
c1x@a��$I�+3AϏq�ځo�z��Oy�\�:��@�ژ���
 0����mG�1���"S7����x�],єA �W��3�f�a�xA�j�0yB��k�^������2�V�x�	]�����
��`�+�� _��E8��&�΄��-\��+������S$�l��d�t#�
F]�^�k��	!�X[�V&�[�PwJ�vCc��D�o5r������]P~��cd��\Ei�}��.�G�
�D�c�~A�gD�����^�X�r��~N�k0�M�KH��o��"1��iIĥ8�P��P��'\���z���Y����/�A?_�*�6jg�l����Z~���>J��0��҄{�����A��r�E
��������;u�kR�b��c�r}�8债"h3��|�դ�r��⢦�z�:����PU�6_t4q�sҫ����!LSt��+��#�Z���� �������_�;U���!T}�ϸ�2�,�R!?�0���M��<w���³T瀋�.���Ҭ�QC�6g����|��h�F�gSs3P��G��e��e���AD��e�х��%XV�tq��̑�n]���o:._�tw�X鍛ԏ��9���I_��-��#�}�Fk4��F2����m���N�p�����F�\��_���3�;�vF<$�8z�*��K�$�����?`l�\�`R�nn�t�zY�4��aN@��B�r㬵�j5ƪ,�Z�_+�a��{�s�N='�c�gE��F�mKH�sٴL�6��.�rO�pO[�D.�J����-+t]�K�χ�k[ny[�
�߷}#�+RX�C@[�Q��+%�Рy&�
2�8d��и0ʢ���k���Ȁ���k�g��=������������ D����_jIC�all,g�����t8�.M�&+j����1G�8�������- 3j���@�/;7�=s�)~N�6-�5!�)h�e�2*t��%��!pZ٬
�����/�ggo��=�x��/�k��X̴�zܐ�>���m{N�K0�RI�IaN<Q�GxB�W��r�W]sK	�3��G�#�.����oA���G�$�:-x�v�o 9��Te��rb��R�n�
�d��aQZ�ܬ�(�1�/s갼S'hޏ�.T=�g+��8���"?P�r�2$�C�[Oŭe!a�X5&���>c�ﯟ�+�/�p�;��,�?:H�$yN��a�/��T�]:�>�,���\·�'�ͩ>N��?��#c��W.�*Av-�"Zw��r-f�J+�|$���+�0Ƴ����g����� 
#��/�/���.��E���G�i��A���.8;7*ܕ�6|�[J�-:��7����y0{͒�@ >K�/7b�uC�c�d✪�w�6o��L�m�/ �~�K:��.4'i�}.���Ѻt�Vn�S5ΉY��QZ�؟��+��eT���K�+����$7���l������L��I\[@i��. �ʝ��DX�E����p�}��|;k�E͢�G��h[I�\
329��n
���BQ�u7����Y� p�t�@7cz�3Z곱���/߹ �HC�e�������g��w�y���a+ECqDckݜȈ#w8k��hv!gS��t,�v�Um 0x��i&�zt��?.��g�f��%Z�f8�� �s0���Si�3�k⁮��6�$����LQBr���+_�H�[22��6��Ƿ�YǀмЮP���ۉ/�J���7j�{�����T����_����tns��I ����Ι���P
������?�>s��Ü�H�@`m{��V��y�.�q����ݵ�OՃ؏ak��
���G.�o�>��3.jڶ�R�i���R��3'�(�q��?����06��ܭw���_w�@Z�(�Ơ�J�5�-[N��]���9����R+���Y�ݠ�q&w ��׭�q���_�🞣oӈz~��͏�!�]���2�X���n+M�VZ�O+f����m�-']��:&Dq�>�����Gf��L��N%�O�G��< �g[ ��h����) #�����E.�Pu+�*���3<|�Ku)i�����m��Q��Zv6;��{�	��o����֝@�w�F��cu�
�d6?1���WX��]��PM�M�L]�j>S�v%�(D���3v4�s�`� �Yկ ���99Buf�E��i���i���]�h
 ��i)�"Q<]�R����7�|�M�Y�;���C
�Am���zDB�1[��#���z匚�gs�������b@D��BC(K䑍��h�~~�н̝!+ ��[�fĀl����(��#[>���lq�<V��-< ��-Gq+�*&���a�Wmw���P;2?��-��� 7��e�Xg��/6ט	O
m>�����;����X��@ �y����[ ��v�^iJ�kPh�����U]<��K�08V�tm~,m+~I��f������Y:.���R����P�����f��h�WQ�S[��+ Ͷ+$8�v�S��l���%��V�%���ԝ�1!l�m�d3���ȇ�2F9嫶ߦ�5>S�y9?Il�O�%�KX�C�w�3����4x]�V D|����e�Ur���~sN�CBl�ɼt����Ʋ��t��^��B�Xƶ�)�z��K ��� ����Q/�+��S4�w��R[�����b'��,�5mb����W�^��p�A�C�eU�S^0�w�Y���;2e������\��2�6x�_����#�QY����v�����x�`Qq�.�̕��55J�=@�{{���B��'��'ߦ9��I�+ilO�I�'S%?� ��7�S>V�zU ��*��Ƌ�wt��u��$�$��g���J��}}�]�G\���Ñ���O�~Z^�"繨o��;�;C���I�2�+��@�R�8n`�N��Mſ��Ys|�2��t'��5W�M7.^�w�G��Y�eD�A��K��f�>{'�e�8�������g��ϡG~�����\�N/��	��{���v�-r���`a�y�����$k���e��z<�&������;�K;�rv�2��z��=�
�$����7�j
�C��*_�y�>�\�ӆ��$���疕z=�j���}�^ȉ�����3^�\������t^V!>�S/��0m�/�����e��LX� 03pd/]~���(���Pv�ɮ.�����|�9��S��j���]�(�J�{+ES�߀6��i4u�zw�+��^�"j�� ������:����[�:祦�E�z�6�����u���m�]�
 �y�,��Q��=�Ӗ�����R���EL��e�?l�#��{�PK   ��dX�Yҙ<  �<  /   images/4c2bed1b-fdcd-48c8-974c-5402e9db5193.png�<kÉPNG

   IHDR   d   d   p�T   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  <!IDATx��}w�dWv��UΡ�:�0�yI.�rI�r��ޕ	� �0��d�0`}ې-@kٖað-ö��,K�Kr��rH�p�L�T�Օs��s�}��:M���B���(N�����{�=��g�����_�wԳ�y�~��,a���~Vp����L�/Я���ߔ����[�Z��F���i�A�]E�/�Ϫx�q��$d����9}�޵E�����vL4�t�1~�F���-tm9����}@�{�����׽ �C;���f.Z�=*M��vG�`��?�{��L4$��rf
���p��-�˗"6��Z�Q���s-��,�ZԆZ�A��A�U���X�A����6����{���j�����pi8O�/�8Emr۩���� p�M�3���V��k�6�[�Ű�S���3��W��r[�Q�>�vL�5�Gp|B��G�Y��T�'����Q��m��*�q�g�T'A��o���}�����3-�*u�p��/��X��x��p~��	F_M��R�Hi��F��/��"�,�����;�	ahwY&�Y�/9+�\��/ML@6�r�_rN�/E�q���y{���99���ߊZa�Z׋bx q�S�<�����,][�mj�����AdBQA�cz��4�=>�d�����y<� 
��LS���+Vض�1�vӄb�&�Y[��آ>f��>:�E���ȅ��x�@�I�c���h�l��Ѿ>$C}���n��I����������<�?��@ QB֙�6
�2~ud��������y�"�������fKV�qD�E�Pg��H�5O_w�V�k���Nr�@ա{�Ӗ:�;,�v�ф��5߷X�:�wm��"?Վn���)�>�t�J}�4.��߳ji�aֱA�IRG�a�Վ���Zm�V�)]�;�ٗ����4�w&ۇ"�a��;kxs~/�J����獏H��zWdp��K-�wzqj�,^!��^m�)��A�(���&rDu����Ď�Οo;�E��Euʭ������\�Lu�6|y��f.l���F"�����N�d��%�5u�i�}�T��O���Sm|}d1B�Q"8&����		��6�����c'�D}��h�A��L��ß;� V�/L��M��C�'|h����~�����O��b��M��:"C5�E�E��&�:|�0VM����}��c�0BB��[+xoi�Hd2�����ӊo���*��m4��S��hB���'"n+�/��X��6�r�p"�ǫ�YhyjS��̠�rߥ�&K�.���VSV/`�ӗ��_)��W���K��mu7��T+�x��k�٣�0l����?�1�A���!"NHiR'.'�\�����c�yKۀ�H��XS���]B��"� �zCd��qd�"�J�����`gR4�h�i�����j��}^7�=2���Aa�nR&�v�P�V���]]�іz���ֱ[Z��a�t�M�wGS$	�0��H=/)4L�~��dk��E���N�	��[�������;=���iK��N9|���pS��W�]{�w9{����TS2��gJ^�I�US��Y�c���Q���ȟ�������.�Nw1G�*�Y-n!�q�|P���P�������<���U&Tv�n�bE%8 zH9!?M�PǾB�K�[��,]ߍ'f]Ң=�3`�ֿ�`n�:>�߀���h�wZ���ާ�ͳ_B��ƓF0�o�?�&��;����,
��7�75��b�^��p���B�; ���!���x&�Κ	lBx�6Q�Ҕ��@�RjuڤN[4)..����A�vh�VU����j��ʤ�N�}����c
�٤g+��mq;O:���Q�d�*�4ư��#���Ū.�
Q�Cf�N�Sx��d���i\����͜ �̉0�}A��E������Ӹ�q[ɢ��g#�=x�x0`��OO���d+rﱇ����]\�v#a'�}r����B�&�����q��s�x��E4�$��4~��1�mVp�NB������!���Ee��[7Ǔ!_?7�Q`�4�[�N�	�-��˗Ep�k�Up�N
�b]�����v��n4;4�$ʕ�aGh��˴j�Ɗ�P�wp���jJk�w�7�b������n�N�$j��z���n�'���	a-,g�~S�����RG�����h�p'�ɜ`;���l䊢y4:wsx^Ԓ�qg)k,}z"Y���t� ���bVf։%��ŨS��q{!���F���N�Bu��U�v����dCdsY�w47�y���+�o ��K��(G#�pe3)�v2�Ù�Ag�tu��h�O��@I����{��[o���=׎�s�T��ݷz���s�r<�['c�<d��y�y��$W������JǊ{�Z<�N��N��'�[D�����Q?\.'��R��bnz �k9��J���و23�6��1K��<��*zL�sS!"$+kY�^��A�iE��ŵ�k����140ؖ.���\�VD�VwIp0u����B����C�����`s�ŅP�H�7p�<�Y��W�w6W���}6D#>���Ա��3:�%�^F�T�:!�b�+����DnT*�p�W�iXv�@�ae=�Z�>����06��i�[2�~� k�(�2�R�;�"[�.G��Q��_i�+�@�i��z�Hȱ�^e:�NXe���E���^���Ԃ*�6^{{E�<���,�M�+g��^}k��N�O���K°�s�&^}sYد�	�&=�+aI�ۨ��p���k#^�f|Eչ�n���H:K"��ݠ1�����C{`c��{y*/��1)�������t�~�t���>��ڒNꪨ�������~��p|����/�j(^;�B�*��}�)�}�kV����BuJ��9�1?s� ���u�g�#���N�laf|������˖�#D��Z�Q�G�T����@�,�p.J!���*��Z,G�վ�����"�F ~Ps�:�tw�o�`ǹv7m�Y�~W >sEX�}��?U�0����3O�!��2Q���=����t���X��������rWo/SN��J���?��%��/�p���g�Ѩ,��3j?��"L�&�*��ꝝ:{Y\���+N<��6u�?�߽m�.i�s�~;wi�xp��1�oӏ����:Q����V��Ҩ���!6� "�e�2qQ��GN�M���5�EQD�:��͛p���n;�FϢ��zؖ69�6�v�j��'6����B(�,�~v`
%_c+W`ir�~�� �dx�[J>��7Lv���5�����mhd]n����n�T%4���,Fׯ�^)@'�=F�z*Y����\t��QtZF��N8��@j]����Pu0�|Z���7���9l��]HJ}������~��c"�w�ц]A�P%�{1[�p�6�J��F�2��`i7��pbЉ\��J-�'�,Y��ln�^�`4��)���y`�����q�?��|���I���H ��f�r'�:�M���P��a�G$��ڦ�7���ܐ���Z�ҙ/��p�j��ULl^�Y�t	���('�E8�6�nl�E�ϯb���q��!$������VR({B���L�^�܀�r�+ET]~�hm#ra��ۈ`�k�� �,¶Z�ꤣ�˂��-!�
�� ���G���0��8�
M���C8B@��`c��PfvK�����\�9�95tn � |��U��v�9;�l�G9��ӎ�H-Z�YZ9^���b�&ןۂ��j��4���ؼ���Vdx�3SBX�*R�pX;���^߄#^��Ԣ�H�Z���I\���a|��:<��v�8�%b\��w;[�~�rf��B*��f*G���� �62��2�'OObiu��"��2�s}�`5���k2֋��l+��c��Zd�᪕D9���N�݁�慃]�7I����DM#g�7byēe4�:G��n�𓷗TΔU%ܸ�W����R��6����"E��GD-�zQz�ݮ�7��l{�:�Q[�\XU1fk���F����A�;M�����$��bu�BmLm����gu�~���.\Lt�^�K��c�Mr>o��4�%r:���r�YU���ҁ
پq~Y��9��ŕ4Vֳ⊇�J���W�0���ܸt5&ĭ��;U�Q����S����D��_�v���<��VH����cP�Q�؊ʇ�h �|��9|��%ӷĝr~�R_tl�J�=�g�-�FU�i����-6��I���N��_�6ͩ�M�2I��\⁤#�k��x�f�F\�ۯ��[�֣�B��T��2�il�o�y�X�Ҧ���� ��W�o��9���|�{���o����!>YO�G��iS���%�9n��v�fh��{l�3�z�����UܛW��C�0�e4b%�
�;3��e�҄.��)Bm�M����YU���ÁvJ��a�hS��~M���t��;׵�TL������jL�ŨO��h��a���Wb��،~;�=ZT��fv��h,��~�ߍNw|t|�Z�7�B�c#A�>ś�W��_~~7�ı�Q��������v�'�G��g&p��
r�<v>?3��W�f8��SON������@����Lb;�ǧ�s����\��]E�����_����1��j	�<;7��,J��a�K/����M�n���'��V�{��`Ѕ�#8W�,�~�{z�L��H��D���bjS��s�ĢR��TB�V��t�^��ޚ��$�2�ˮ�dKRO?O��f�����r�X�n���=I�؋A��W��n��P��Pˊ�U�1u�o����L�Q*[�T�Kv~9�Z�-IdyB�<	�<iD~��-q�1p�VcG%��J
B��:T'/��wUS�Ej����;u�)��l��k��-��R���r��f�PB Ğ.կZ,����G��I>���i�B�;�,)b�fdQ��K�b��Oi���	�n�_��O���/�,��E���V�����U�g6SC*�Pqe��O�5��gRy�(b ��m5��ZJ7n�%�Y�e�a���˕n��@�]9�x���[U�\&[E*S���n�9�%��TuI;�������wR*�N��F}o�2)Ɇ�P�6\ү�e��W�c�����ڰt{1���;�I�+H�U�fU)B7v�K�>)Bܯ� �0{�K��x��F���;�7���'wN0ӏ�����=��=?�����n��G8�����~��~��~{kSIZ�����W#$����2� ���D<4Q��j�
`i%C�TE�N����o
�c�|vamLU,��L�cc#�2�YZ���a�!^-�n&&�$�{0�3��olW��Cn�{�=�~���o2U�VIE�E�NƦ�J���'6U@�����a�)�@Y^�K�ˎ鉐����.��H&�i��dC��l���D���<5%6YE<Uy9�t	\0�=q"�8���J�	�⣑��95<�e����	BH� �c�x��d��Uz�&���D�*-ݜ.��Q/	L�Ĵ�u9	!ӓAl��Tu�H�>:>��Ԝ>�!���ؤ��V�A�i2s�H�l�P�E���L������R&TR���QѸR"���|�&�����M�.I��G��ŉp�%M������a�1A6��Ԩ���8!p��X�&!�d�,��ki3��\��v	b���p�d�����n����t3)��w���X[� �Du��1���7�ƛ�2���)4.ܼuEVN�����c�.��^����F�Կw7Q$�i�'mj~����!86�B��}oI`(�ǐ�³r�Xu͎u�wt�:^c^6��N�F���RY���!䶽�	=��>+�p���5w c���!�� �u|�
	�waI�CC�yC�B�p�}}(����;��|tJ,n��'XY!������$0.�XT�ɑ`��駷���Q��חu B�x��� ��a�8�<��Ut�N����Q)��Q�G��Yv��ӦӃ�'����֨�u�2�!�h%�$7i��N<[�.�͒�XB�XQdJeҤ4�����e�[s�କD;*SL�k���:<X�>���l+�8��O%T7]>q�>�ؚ5�L�fCH�M��U=A���"��^Vf�@�������ɺg8�_�v��O�p>-��VS�E�t.����w�?B` ����'���ʲ�5��tm�C���M����fO��r��.R�`�����<
��ڦf�����'H�hb����~��#'g�mQ��1�s�䌬V�V�j���&b����􄔙<LMMI�L�۩�����V
�����#��5��(7#��f%|z���w���ԩ1I�mV�����7i�V���cjt\��4�fT��\��-˶���;4�Ԝ)W�Ht�V��o�a�Ӣ���^���3���[�U�F�������rЭ\Qآ��fr����좡k�ɕ-U$A�ZKU�5�����X��\��1ר�V��Ѝb�*2�"m %�2������\"��D�s������Ɛ+�v�#Cv�Jk�p4�2���
YJ�>m(��B��
Q���g1��Ƞ�M-V#�'��������*sQ=�P�Ւ�攫CS׬������-������-T�����c�ͅ��{��������7�ĬRn�H+t���h��5�k�|h�R�1�Y����d���Ų��Vi^���n��Z���X���A���
U������B�6�Y4Ͱ��}�3e
���1)��Rs�q��?�X�����>lV��l����g�t��s:0��Z,%��!�!�v����r�pf��#��"�������(��6r���Ǵ�%�@/�e_�E&��!%'�.�#^7��
$#^ɮ�$����G�Αx�TR�r�E��F��E�a[�v�v�.BX�xp��͌�F�)�$x�0B~r{ӑ��Ju���q��ۅ��7�L�a�):x��e+?�r�L�\Mij�d���'�[x��Y����h'�d�uy��͍�=0��$il���-=0��O�������>[E�t7�줕;��-��N���7&Rv ��x�F����Gp��G��-��_�\���t��n���
	9��ۚ�`M�7�0�3��R�[iYE���y�
V#'��"TY��Z]� \�g/��x�,�/m�������u����am7�g���l�@�U��-v����]��L!̂~pmI4�qZI�v_X�	Y��I�Q#7iaU�����k{k~]�1U0;b����k��O�B��oq1�%����O��խn|��^ib[|�����sA?� J���\�t�glup��`bÛ7 � �2 �}	-�+�s~#�������t�ڠ�=�uD]�	ZM��P�d`��gdG0�P*#�4^!��`���1ɶ]0ś*0?�v���N�k��!�_Tj��.�SMu�s?6�gfa��MFˇ�.�Cl}����5�1��*	c~a[��N�~��ܣ-��܆�g��@=z���S+��?h2{���mjn�C�֊�|�/���ae}R��;FF|X^�vm�.Bx���b��F�J��Kl��e-�(G�����3�BZ�N���.c+�"��_�zekY��ph��`�
�B>���1�4QT�7���O'Um�s��Ϲ���ە�Э�����b�hyܨ��*�bV� �	[��$x�$�WHem��S��f}*��
g����[����#����i��n{ �j�Ē��|tB���+��5hs��Y���p����ʥ�ۥ�8]4�>Rt�� �f��$�g=��c�]?�9~f#��o+��X�_؆[o�N�l�䇫V��]Z��滚��q�W�02Hr��X�1��)N�)�h\ߌ�Q+b,���A/��!vP'�-I�[[ɠD���l��σ��:թ#���L�YΪ\Vy:s�"Q�뫛��C��R� &���2L�r���:��QS�1�_3�6s�T=��ņ�k� �&2��s�F#�><��8^y}^�y��9�I������aHN�p�r;�?`�����U�<��0������{��$����iU�M�qz.��d��Y���Gp��<�*ms�q����ĆP�J����bm͊ ���|���r �q"]m�C?vKxH/��޵�i5��h���y_���Z����ʹ(
i�t>Z��b�?�Ӏ�c��MRm��$0�D���l���b�'��J�FZ���i��j�"�(�)�jq:)����˽i�=�26q�J��ӊ�5.�FU�:���S+-��F'U����4�S(tm�C�z�!�`����h`ff�dzU�A2��G1��\��ᕨ&���A���kd��`7v�r�V����l�Ri)�
�S.����U�o~��즱r�7��mrUVPذdYh��''��R�o�&V�^?22"�R)"�"����
�I����#"c�����G��ȥT���Q9K���hY��v {c%E�b�S��.JEޅsoH�c��W}'�wDq�%�������I�lN,3����K:�C����Z][��4ٓnn>��e��F��n�v���E�����/�o8��G��xkERZW���x065-	ܙBE��#�Ė����� F&�d�K*�����T��ّ�L���K,q���O!���s����:��"j.�n�����nvM����,�xc��n����'��JL�fϝ���q�bL4��ω���װ]P�|�j�v���H���h��Bx�U�p]�l����݊c%VBy��a���?ڔ�-F���f7�v8q9��d�J��Ɂ�~�ڳur�sbtѾ0�LDnZ�=������iu��>�ﲻ���F+���.I�j�it���B���L+��*\������ժ���!��o$�]��DI���E����l媵0�����q	���d�A�R��>�dm#�UQ��Z��u�E�^2Uޗ�����)�L�u"�� <��o��vv`��'�UI��5gnz����|�������dҐxW��cW�͆!ː��`ð��`;���L\V[�X��k���I*g!;Y(fI��\��c����}\��MII�����ϫ�1S�5q�fJ�u�T~���N:)��2IݔtRbU,S��Ji�
��y�w�٭1��]�Ep��;|�;#�wlGԱ�JtI�����ݲ�e"����V�3͔��X2!��X���,?.��>��h`1��{��M�Q8=Λe���K�< '��D����ٹ��#*m7ǩ�*L��#1��+��+�܉��J5��q�m������+y��!�)8��eki�$N�:�?>M���ښ,�[�1��mv�Y=@v�s��BI6��I�څ����i��xDvh�*�sf�O��8���x�n�G=�r�2��'�#�ƚ.(eal( i��Y��^�nt�Sa��a� Y�|��˪-4;]v{��M��0<K�9��ύF��!�:��XečGūo,v�e!�Y����Oq��<~��	�I�u��4R�����������4|J�&��SD	l�����03<��o�m���"u��L�$!H�є��T&OF^Y�F_�EH
`m=#"�.~�Z� �WH�ͣln�e��Rာzf�l���2I�5dN��-v���a7��q6���ggGa'byg%�B՜�|���x��q��%E�λ��K��ۋD�-��슇<��x��'�D1������"��'�q��)��7��h(�����C9	��b��jG~`7n�*���1�0l�����Eۚx�b
￯�I��!d���^�D�����?���u#]����i�����2�<,�N��Iy�b��9�#�h4�k^͜���z]	��	��ۊ&�wXj���|�!�z,C����ΨY���IM�Bufe��X)n�S#���F��2Y��9��^�z+��0��l���dU���矗l�D�~W�n�`�b6�>��G��$��F��
{���I�ȆG��˔q^m������o�%�ɮһ���rP�kђ|Q���@���"��A	<������*�{&N�v>��&���0|u��2U�'Rw��O+�����v��'�?^�� 6BeR8�Cn�m�j�,�����vՊ����Ѷ4����$8v���iV��b*�|U��QR�bKH$Na(�q��/�8�vxZV�N2���~ߣC��H������Y.Wd0��q��'��"����m��9�{xJ~�JZ��e-�g�剺��R	T�'�䭷�*�]j[�$���a������vf�C�/#����_�"�k����v����� �!_ؾ�p���0�:��Z���@�`��+0:�Źs#x��%!Nv����Y�V�{N��a�Lk2
+���>�K�4b��Ȝ��7�i�J��Kg�D5Ζk�x�,��d�)@�.U� *�Շf�B'?|�^��ώ�q���e��o����,n�ra���ĠLһb�V�J��DF�3�ΐZ]���R��U�����٨l���kb���������*�����sC��9��;Kr����iRl�8�y�ռYB�9�'[��J���._׾D9��Q�Β�)[Wi��x��sУ��n��n�B��-��/�=�ȩ0���1�1S>�ʼ�S�����.���E`D��5|�N�a���b��W�BP�>df������1YyVY��&�|���c!6ʹ��.��fsK��Z��9�q���e�=��2SmY�=��S��n�KM�!��`ĤHf���4y�	5��e
��_/����į}���B�y�4�����'�[��I��"�W��5��8Dlr5��Y���Fvݨ|�F��W��E�#���+T���:��t%.wx\�3��{�3I��dF7G��i�����4ё��z�YlWI�8I��F�&�?��AA��2�T������9!c���Ē�8D�&+�$tRuyųO�3L:����m���+��q��9;�^~�e8�nd[�<
cbr��|�r��{
�(ꑿv��G�7'}�3�a�;{����S� '��bG��tdb�u�o|_�����ra}�R\����	zq};'��sqy}]Vq`xL��lv(��G���?� �!�
ae%-�a#��jx�ױ�O<���	��-"�G��ժ��_�9Ƈqn�t�������x�. bq��ƫ������+Ð�E�i}	ډӖ���90;��fnw�	7�����_�u4h��>d��_t��lq�7���'���O:�������s����dO=����ΝU��.2BD(+�D��V�'K�۪ֆ��] �������h�4��f�M�E��_dIa��}欘�]�[޶�}p��TY[5��\�]���;���z�Ñ�G���]_i+��;w�嵔������+�iUپ	d��#�Bj�`t�3��H��Yݣe_�8��bU���:����P.1�_��'�kF��3�3���]T��.HvH���N���ǻ��[�pys{�f�E�ʽ�q�f�����-���o~���o|�{���S�ҿ�#,��wمۓG{X9�>�oob�^CP���x�����l�c���p���b��{ٳ�r�{�=A+e��� T�'�K3��{�j9n��o>yn�=�����i���f���m�#陏���� >�����J֪���/�d���_"cݜ���a���D�nq�����8�l�j�]W
����=:6�]I�j]�1{V� �����w/{y^�C͒觩���_�?,�n�G��Kcu��0�sш��8�R��*�[x�k��6\���xr�#��O��2B�[��oa`0 �|񉤎NS�
Ul�o A�t黝� ��RoInOW�Y���G}��lww�Z�3x�}�gB��!�]X���&�q4�����:N���R�.��_vr��BDl]�W�Ӥ��X{�v��1\���甛��;k��� ������D���I���)��);]m�d�?<�/����-l����l0��܉(�Et���5�:5���[��8NaD���a$K�|�Z9h㎜�P�
��!�'Ǉ%�za9&�k��p[��^�����}NSb43ys(���+��mލ�u�#���˒p�V8�F>\��W�ز����q����.�¯����E����v{_��?�7����ߒ�h���X67�'B7(�a;U��8v\>����x{A��l.@;�D䦾1����qX\C�S;R�+��?��XŊ�Dd�v���7�h��7݇|a!�֟����1����)��~�]��ϻ�yryҘ2Bk�O��/�1x�fē���1��4殜t��0�p_\�a�p]^�6S4�W�	��e�w�gm������k��~J�]�1�KG]�X�37'��6��y�	G��49�����һ~�*2���''i��I	�n������[���-q�������a�3�������h��ze������1���b����d3��ͭ[���cdX���OM��!8��g$J�k|P`��zx���)���=ލ<L}����l
�}��9��7��N��H��F���pXwe6�W��+QNk���ĖfE�; ӫ����=t��0-=G�ޭ��i~�%�M12�j��7Qh��7�D�7E�55�'��9hŬ�J,)���4C�a��U�����e#Db����{���f���[ż۲�Wm�S#g����w�$��%lI��.�p5��~ �pa9.D#�E��R:�}����߷�hc� 쮒�jF9.Q�tI݄�3���qt8�-d�G�S�4��-��v��Zw���I!-��W�%��bQ�L�#��H����DV�ov��m]��)Qv[�IwY�l�4&��F]���n�M���y�#�n~���t=�>�m��#�6��R�p���:��3o����)LAߦ����!\�|1�LkG�wrn�S��	�

-'�s��$�5��cEDس9[߆g�q<����!�ye�k���~�߆�<��&��r[��~u���J��Z��׆8��q�|o����J�*q�?�n#Q���1���1i�?J��P��oD,�t�N����'���_	Q�5�q�j�>hÐ]��4mogZx&lŋA���?J��~����x=G+#��}6< b�}7�$����8wXǏ3��b۔���k��`�a�}���2�Np�.���i/�
�w�K�ة/�(���m�kM|P�Ddב(a��������]sjv�|F����x{���x����[�xdf׽^<�!�e�|ix�Q<f)a��>?7Gu\x��X��<����Ƨ���X����N��M�_�:����{<x12��kt�ֲbi��F��,�B_(��ãr@�x-����t�4��V|9�#1�Q<��,n!������lX񒿍�;�052�GQD���
E|}�nU4Z��V�Sׯ�s%�<b��Lf�٦�g~��c�y�.�H���х���p�Շjt\V��R� �I��YU"��Ն��/�2]�Z�x�%����^��p݊�F}^�Tl(u8�
�IRj�L����v7h퇝�B�C�����-�r[Ҏ�*�WM��v��E�Cͅ��ҽ*�B>���r�ÉR�Ȗ�'7��	~厦�#o�a/2d��U�Ə����xUXSc�Z&�Hj��j�*6W����P#!�w����v�ŮQ�a�����E��O�V<:H+���Z��<~���$+�&���v<@u^϶��񽤎�"����z�)�=�'f�
��mҽ�l[��1&�z=�;/Y�jaL�z�f=MY�A"��h �-��q�Bd
���UJ��/���0�&V��:)������z�%}9"$B��ݔ�A���u6>�$Wm��.�������֦0�H�G�^�[	���햮f�c��˥ӛ���NZ�����rKB����}7�V{�5���"Ʌ�̿�Ziz��4�rf"#��콂����|����)��?��H�Mۯ�0A�Ih����:�g�}$�݊U2����*�����(��8��Fuj4q��<+�{�O��4	��|�3��*^�P�A�����A�1����Y&����
�-5�^��QI��'�:ت�����=.x�i��1K�:�
��ɇO4e���h';� �+�n�k��z��X�1����%ٛU�
�σ��is������Pm��3<�O�����kr� U���c0�k�� ��aA�ΔӖFJ�^x�|
���-b#t��Y���{ۚ��6_iˎ$_�,_z.��(ٽT�F�UR\MN�	tjď�(P>�]/#����D��J-kX�{���>�4�R���氪���;�A��i��p�Y��:����<�~�|8�||A�B]�^�JY���,�<�ejO�`�Ғ��Zt9&Ր��{j.��̈́��˨4
�|o\/��h
%bq���"��a��w²�� �%�ɾ .��ʟ�a���ύ��8q�������<1�W�Z�Vm�$=��4��S�����(�TgI6��6���,>���B�.�p��Q��_=t/9�S�^3�*���8>��W��Ŗ�Y��n�Nz���ϏK�i����zWn���Y�oj>;�#�}��L�����W;�RrԒ�� Q#�~�T��lF6A�'!Z^kVY����1u�g4'ǋw���ַl&�,���7ն/t$!/�)���Ѩ�lq�Q]\��I�?k�id3<x���M6�{�/ɪ�kb�z�v\���Lao�{�?�	gO��/'�8@ƙ�ʅ�6d���|�D}��Q��|�����f��N�|��2�+��_!���X���ZVG��M|�U���KE�$
���p);�
QP�ừ��,�����]5�Ă����!�t�V�#�2��2`��g�$*E��Qm �&ɚ4�s�m�Nu�go��d	ir�6�T1%ؙp�@u\%��C�uw���j�;������1K�|]�/8g���#�_X�������a�W!j`7#�J*���>YJu#dJ�O ]����@?�޲�H���d�F� ��wH����K&�\hd�;���M�9�#�]�J7= \9���=!���3|{d�~�d�5q��˖cJC0�q��h%Z�vҿ;����"��.�O�v�ٛs@��>m�)7��=�������0�-����9��V��    IEND�B`�PK   ��dXv��� f~ /   images/4d249bba-3190-4770-b321-fb8fc027a237.pngl�	XS��=��-��P��(We�@�U���2)a�)2�\�N�'"��@9P0̓��0V� �� B � ��oZ�����<}�޳�~ǵֻω׎�Yl�z��[1��9HH�TKHl	�,�䧙�g�|�+��f�O�f�����ly:TBB�9�練�'�*�9��F8�-A t��C=�{���f��A�ۡ����辱Â����{N���N������-Ү�7�g���װ��6���������7!AAQ�}�C�����w4����K_��������R�{�����j1���}{k�<��=1�VF^x�/8o��P�p�[L,��^Fi���0UX�����W�C�ʰ�e9�N��'�"�1����J3�����B���Y���@�ڌ6Fն|/e���YMFb���7Q��yp2&�(�0�6��j����Հ���_ڟF�Ǡ�����c�t��ZD<$����}��p=�bu�l1|�m�)L�N�Z�ش=�Qm_}* �5�)�6�dK�.�
�}s[\�g���L�
Gwj��Yb�>�T�n"X����m�Er�$	F6��fw�oV�`r�������AU��b9��X��E;Y�{��x�nް�m��C�qF��p�8ƽWW��^�tO{���1����?
�1�*b�~��wң�(VN�[���i{������ ��91��\�-~�sA8�O
���R�x��BL�ġGgº���j�� <��qx�V�{沴1��tfo��qҀ�aHW��@p��H��׳����*x�
&Έ��X2����]��;_�O6���P�Z��D_;j�g�9f�몫�fQ�̩��22s��ܾ`_�?���0H;�Y�\�ЮB� W�?G<�-
�ѫ�С'�$K�<�lɠ'�����D^��@�P>�p��9۸�妡��(�n�O^hb�^�a��:�*��GA�0~���A�̨��r/����
� ��T���R�>�z�
��2��7G�jL(�PL-y���J�#ݖ0|6\�ѝɒL
��/�=����FZT�GA�`���[�8-���P����B(���0��+:���%��<XǞ��F��ʤ֜�����t+�&<у�R��(l8r�9��~�[���@r��2�4Qs[������^J�+��s�
P�L�|�H�$t����Gl�5wZ���v�]7�௠�2����'��|n��K�NcB�������œ�=�O��7x��̹v	]�+��6�ryS���i(f�=a!Yx��b�;�퀖3Qk:�����m
c��AV��/gG�,��WQ�e��^
(��WupA,��}F�o��5�()�75�t��r�U�eo<I<�s7/��a؍;:�-�J��c&��>��:� �H�ys��q�5�oO��Q�E�1�h��h��~���p���/Lg48'�����yb��J���;�70�����Є�8�)��G"w�\���*��á�|<�1��Oq���5N�7��3N�	M�	�x��wJA�I�AS�_{�ǰX�4f"&-�nӒ��Wh7q�>�\,�z?�Ҍ���:�
���M({,\���-��\���ip������R+np�4ބ��������
��(�Tj	O�D��0���.FAÖ!X| ��(|�cA/x¸�bt(7��$v�'@���d� IܑUYZ�<E�F׬|�5~_�j��l�$��p��l L2�$��M���U�#܇�Z l;O�aV�\�e�p��8v�*.�-ʜO�%�t	��bA�3M��s7A=�	*e�&*�d��c��P�s�4��w � ZJ���2p�$v��ʵ/�'��QP�N���y�r�S�$��6�(�{��)�Ѣ|�1 ��"ju�౓؆�)��q��	��!�fd<>�B,�#5{�'��}S�;��d���B�x��~*���۲4�*��%�ݟ��0puEb-�����}����,!Ḡ���3jA�X@�{��9ǰkA��_u���C���Uv������8����^b��`���Z[{{NFN�����fR��M��A"
<p��O�̬Q���@7g�C����L*/���g�Ν;o���<�x���ӧޣ������fM�7�.w��$��x�p�G���e�\i�T��=��-��L����Km��*���'��m��t��Nc-�O���0V"���&����������Wd�nl����j/�~�����Y 02�s��]*����E?�'CY:ї�)�//'�������K*舃��mɮu3팆�t9��\R1Qy�nv󐁢�*p{�>���=J:��a�o�S�ʽ(���#0.� �-�����F��赶�֯i\L��h6���Nt*�*#3��H��ȵ���>F]PLla��a���㞞}u�#M��ȸ������ᄞ�R5^���[<���ZҴ�Uߕ{wt��dge��v;��� �ȋ�/5�LO���I���ynO@{?�.�,�A~6u0G|�a��P�=q��P9h
ix�~��|/uf�Jls����p�%���XGz�ٯ�8��Og��C�ePG�*ãQ/8��z���0�C��>��7��6Ӏ�97>��&���%�j(q�A`L��<	k��L1]`�����}=�R g}yᖸ��J�=��� i�A�탢��^#{ל�-h@��)7�2�K��W�^e�K�ڔC;�@Q��	ۤ��1����+�NJ�ݎ�yL\>Azس�Z5��k��@z�H� d�,.x=���Q^iS!�F���ȕ����4Ǌ��:xB8�Y��&�&��Zԍ�۲I-)櫋�����<6��
�6�i��W܍��yF��/�N�^TF������=�i��t��|`F�$˟Z�Sf@��t�XY>	*n(lچ�Z*,��C�k`�=�E"L��{6[����S��
B[�~e�*�w���`O�6=�8t�!Sq�����^}������fO��"�I���ΈuHޟͱ�Ep�mS:�#��d�F}|h
��V��o�/�SOF����8���$>���Q���l��N��3#f)'��rCe�9�Q-��s馧`���)&ô㜾�tHE37����wS[�&*�cJm�x�MY��}�cl��7�E�����b�A"]�.��^!��f��d�d�����Qը�2nz{e���-��w�`�s$z�%���E>�qP�w��y����d����`V^�Y�D���œ����˙i����| 7�yy�"h�H0��_
���숙����r�C. X�誀3��$�6Ͼ����R�i�ho�c��m��ZsKQj��I�4T\�$Pv�ހJ�C�r�jζ%��7p�C�<���.�㥧H���f ��AT"��`~�ސ�O�,��Pw����[��6��ͣ�
��(GnW9b�����T_���}�=�������b�� ���ct��2jؒ�����U�cDW�pC����$���c�A�[���ױh7���ⁿ���|k��4�&܄�@y�,��s�*w~�_(+�X�1x��$	~��=�u��aXL���F��;��j��&�I;�oj��ωf�D����\�3U#h��S�s7ܗ?���Eb���(5DaIf;��}opn<D~����D��F�`���s��s.�*M�ܺ�BG_�
aۺBx*nP��ǰ�4kv!z��u@,�(k� 9�/���)�#_�..m����2;w�;�L�uT�?�VL%�<O� �jv�"�J���r�kS��-��X,��a��s��%���s�Gnl�f�]�,�K	R���#� Y��bV#8������ќM�"�L�C)�YX��c��lT[�/(~0�L-�4�96�VP��-Ud�7Rf�9d`��߽@	��+z�_?:�;Mq�� f5DO��$�=b�v��ſ�P��KVA7F�����~��T���2N��~�0PE�F�O�췢6L����<�nw�Vr�S�&W�ϑ���^Pa�Ą�sR�������jf���j�<�p��(�'�4�Q��zZ�c�̿X��F��7[q�U�~@t����w����$r���=�S�=`�. �2���i;W�7N�wD]q�����Tz0
����O�0S6U�KQ��j�KjQ �LP�17�|p#��L�ɏ�@=�����?Pѹ^�� ��b�޻/8�0<uS:E�;Nw%�.�u ��椝�w��3���MI�X��h�L��t�)���i1s]m����F �C��oq�F�9�qh}J&�s`�-P�N��Yw��'��YOM��y�/F��� ?n�KŨ��=[����*-�?M3�+^Jb��$�i�����M��u;��~xJ�`'�o����������a�3���2��R?���������#6'1�"<|�:�%F�`���	�h	Z;VmxC���#rbR��O���4O�3@́֜f)�?O�vm%��Ew�#�����ϑlQ��9�J�&^n�_~����G��$�%���R�N=����H�6.M�Vt�������|������}�#�4%������XC���@���P�뢒�AMӏ�2��<݋sv�⡬�:�f���%߬�� ��*��b�r�N8���7/{��I�8W��r"�3�xܱ���ίw.wH�|��G�m:f�LH1���F�.��]�3�0:�!>ÏZ�ʽ��J*�~8�=�ο�rB�G�}�1��%��uci�v$z���|���ypq$q-t��V�O�րB�v�9���Y�:��>�VyJ�W173[�ĆG�g��YԺ��S�a�
=f�ik�M^��'�\f,�ԟd�Z��	5=ͱ/I���b��8�|:�.(���(��v�E����\��XҶ��ҝA���Q�d�j�D�:2�x�Ǉ/�ƻ���e@�L\�t'�=R��eN?��LX��͉l_f��_��]+δ\��W�Ye�Y�C�-(,4��7-�2u��5Fż��}�%w	e~���# Nt��6.�������NS��wM��:4=K�z�2C�5�Q�_�4��>hl��\\�M� |�2�����U���㙺 	��3�qC����j+Wz��W��F�B�@k�qCC��|��?zX��y�_<l��8X+X���u;���!	��|/�~�ƶmۈ��[C�����)[�ϊ�z���̹��8���KՊ�@5��Q[^8
�\baVH���XQ�a`X��PE�����t��ZrD߇W7̣�ˁ����&2� ��������sZ��.���v����TaHQӈ���,��$�J �zМ�P �ߢ�[�}o�io߾dh������y�����ϰk����N=��a�29J���*�ts l8�(���q����!0;��E�ʁ�ؙʡ����	�I����b���â�~���/E����ViY~
ls��r+�q�ن��  AT��u�"g{m�&�L�?C���H�{��6���j��:���FtB�ٙ��D�|#�fw )�Qmz��8��afp�0&�Gʫ�h�	��ʋ��)�JY��Ճ�΋����[���k���i�����֤�*Fk@�gmA��{0?
�z�� y���K׈���0Ú��68�v���61�C�c~��c*�'�n��y�FK�ݼu+�2��e(��u��3F�nTcO{(P�{��G7gh_��Ϟ�p�O�8z�Dό�	홹]�q��b+#�aڻ�(���k�_
���R*��.���G��~�〴�(��܈����^G(S�n��M%�젩i��˗/��}O���-t_�vm�SO1�>3�عx�"�?�o�4t���u�D�Ak9�KpT46���,�UY��[dj�����kY�mО���TS:s� �Z?9��oP�1r�5���;�ewLw	<l�� ��6�(�x��L�����$aإp�So^N��5Pw��7�Q�������:bL?���D���vgݻw�����o������)� �5#�/�F��|,͍��2
�~�c��d�;�/�w��0E>'Y*͡�i�d��? �k�N�
'���+dj�9�ɽ§��w��a:�@X�j�+U׵��z�
Lz|Y�B^�'4l�eS��M9�l @�@��וz���^l����>�Q��o��B�`w�b���b��2�[2zf���^�L&�\�{����[��d�����aܳ��/��>���쵈�5�S���d_�:�鄧��;:Db�^K���])C� �~_;\���k~
��X��BOZ)���ĜB�6��whWMۖs73�|�Z[�^ ��lfH�L���;��H���tJ�gV~��dV<���~��0�%>�WL���kV��FIw���FO�+�\4��M�{gMF#��cfӑ�S�2���7�^ݺ�@�����"2�Q�'��ǆ[q~�}Ip.�'!��\�<�n
�W(9]1n����&�z#��PB��y_� w����Y�^\S{��}��B��u���=	�̜�{e�cP?��z�k]��B��g3���2�5I��L�\�w
��I�m��|b�Se�Sm�~���O.lB&4ۼ3�sW��B)؂~y}�^�S&�b�΂�RW�;��|�ra]��i��r�k@�OQ`���"�;�I��&�4H���ʔ�_?�]{�L�1gϞ=S��i�����5�)�E��c&��dcgɵư���84J��N���f���Z�+A!��n�|˼#��n��O�<��}TS���YY1�g�.�V� 1� ���N}��D��5J:8�;� F�b,�-**JW}�N�OjQ�]�p#���x3���j$�A�ry��L�������ٗ%�- �f����F�c?+���M���n��:�U�L�	�B,��fJ	Uڌ\/	2����u��bX<�^<��8$�I�:��n�n<n��%֏C�:a��	�O}��%��G.{4zrL����C(��>_x�+��\�%��I���;n|�{\���~v '�Pz��{��޺�۸؊3=����8w�.'XrQ��p&<Յ%W�o/�c<G̢�_5ǂG���+�yV<��C'��[�f��{������h����*U���o�F��`���ͼ򷙼D,V�ň��d9���^�B
͝ȼ&�_�w��	�\/�F,�	�g-�0��}�di #��>�WRW�3��irdw�H��#+�H��/��N܀��R ��b��(�VG�V	I�y�z�{l��K�G�5d�ʟ�_�3��Y����Co�c�zz��o��Qڈ1$x��u#�C�>����t�4�5_�������526!�=HƯY@k�6����';��)�b�,L�il�VwZE��[O�3��g�7v=}�tkϧI
�<n����~G���΀/@[���d��1�ӈ�|�.S�9bs�`qp��O��Z?H��\/���I+ŀ��>��FI�3� ���`���1ڒ�z���`�.ؠR�UC�й��.�+�@�'����	�>��.v#ԸSV�<�q� ���S����uz��X�{��v]O��f�Z���=����%���*��Щ������������e���}��X�O���f \��+U�:WNw�������в��v7�im1��r�CAq���d�ۘ<ώ<{2Ԩ!�w�ͅe��f��ؤ��/�d�K,y��9u�=��hl��G�t�W��|��fϝ��`�k�`�0��A�l=�+v�}�6����'�JmJ��+U��I�q5	r��E΋�z4�*\[w�'}'��m�o��U;.���:i��$����{��'��w@%��q�{1�s�oL,�Q��s~#�s=�� ����}et�Z�Zw��J�?eKa�2���pGlC�}!Y��$��t!�G���a	�))�������\��~~S�7SRxv��wPj��]�V�{/��`�-�o]����H䅶�]	���DZ�f�;E�h�����:>�&����8: �I�c�%��0��0:%C�7��c��Ka�Z�0qY�/y�8b5Q���j~��Z�h'��!7�%��M,�2�簈��������S�]�ČRC"�6NHt�:�Gzr��y���rA���
�C�A�ȈD���,4u�����e��w[�Cw�م	,��}�b�����`rr2S:�����@�;Wp��#r�l��O3Ж�cF��ݔ�x �����֔V�0/cv
뉬[�=K�ӟ��rҨ)�nXM1]kt�燌Mٱ�P|/������j8p��&茺�D�w���6�(�4�9 �f�#�k5��.
���^����j͈8�f�����B��K�̓�=�v�\z�R+���I���v�7��a��-$�^S�b�*}����>�&�E׳2��%�62ed3�0�i�51��i�Ob]�c}?�<���䥘�>���}f�	�}^n�B�n��o@'H��Dq.�������`x^T��@�?���yϦ�E�vj��q/�܋W��Bb=� ��FǞ;�r/��gg
�'��.~I����k?P��LdVN�eB��`��6�R���K�mb�f.	�h_p<ΜȌ�I�p�eJbZ��$���Pkf�0P�K�"�l��n>xY����^��Vi��l���6.f|��Uf�]遗���n����/��͋���0���r���Ϋ�1,�d��{�5�����+��[H�����		)'��/��a����r+C����ġv�"�������}�0���-�)�lKfhU�� ���r�j����	�]�W#!CD��a��ń�l��D*�J�=T������=&P������U��ow��H!�)O��Q�Xm���|o��� $VQ��ޠ��b�Z����/:u�C�!���[�4��^��	��:�mE���7�H=��/���E}3�J.3���;�Y"�^�R(��7����zP����j9G�&'�r�
.5�~��
�������{ٲ1�L'��[ųQ�V0��a�(�0썝�F�ڇ8pT=�/zC�"7�N[���Q��755]���
��{�]�F�ͻbK��۱�0�
���NK%�����IO}mo$��.���R�k���|��LO�����5l�0Z*
����wPN���%n�����g�=e�tP�;�οv��mz�j>�a��bx���W��®�@h��o�&�۱k��SX0��b0Ă�L������������e�5>�7m���d�ơ���>�34Z�Ʉ�r�fҿ��f!&|�Գ�~NNNW �N���0r���<l_����'���b���!Z"�����b#@l6C�OF\�*	�#�c��P���٣��p��K�M�a����]���]�1&6�X��)�-�v�X�6��r��g�]���Q�|:v�>c�'�}5���(w[��-CB�@"�̖[� J��D��j�%�6�kn���a<�/v~�r�ޚ����U8ه� 2I�.Ҿ}�����m �9�b�D<�:/k��/�EwL�!P�|+���A�sJ`)�� �te��);t�frՔ{���xjZ���shttt8�r��xr�v\g����<^�ܰAv�> ��n���7� ��o
��H��mL�ڶ��N�30�����aml�3���u�]��(H���&ƀfkx#���.�Ef����i �Bw�@�?R& �;6�V�<�����%x�����<�M�L���1��w��;�JXn�uA���g���K��Oa;�,��~%��#V͆k	�h��}�\�c:�j`XgJ��D��_�tu����%ڋ+2��ȉ���*�Z@>��Ø��2�h-���1�g 5��_'�jFt����̣	j�<�w�չ��T[�_>����:`��w�~�u����@⯵�;B���FW�8dn����1U���R�/��En���
m*�w]�r���հOnq���?r
����x]���Sߝ���yݬ�nS}j�r\�J�͙��;�C�Y��e$��!��8�$O yݼ	L�F�;����x�ꗒ��z���~��*������+7{x��s�0�?�+���b�<ɭ���2�=T`�F���C?YB��5�¡=�V���Z3���E��׈���&��҇]�j��z���0��R�
YulX�J��!0�H�z��i�O�g������{*m�ּ�M@˟���bʟ|�W�cV`.V|1gOݒ�%�(����3�B�7�U$�C��w����5�Pi�u��
��B;�5i����M�L]ҙ���������������u�@�s���ߤ�@1f�y�����5~�:�'}�탕��F2�KS2?5�$�oO����9C1e���̎�L�����f���O�;��g>3��jD���*:$HQ�yp�;	�IK���5VJ� ��{[��r��_P��d�͘�:���'��d___�4����19(�C�Ńhʩ	�^P1�>/��P���;$y?����1��yq=QԊ�[��=;�lb]��������N��%(��LA�E��Q�J�c�}�i�\+�3��Ä�z��
G�����au�O͒Rl��q[x9�6u��ӽܡ2�Y��]��OR��-]B�5�\��X��7jrU�8<2�hz�BGqv�+Є�{�k�z�\�2��5�ĲC��Y�:g3Me��v��2�,���Ĺ����Kw����H�var�x�!_�7־�Q;^ߏ�-z=�k�L���D�**U�����VZe��<z}d���xzK������cv���MgY���d���\�J�}|N�����~��}w�cφB0co1�	�Y����2cv�Y���K�M��tp������j���I*�n�!!!�D��kmGH�%<�E5�f*���m@���:l��zs{�y����K��0�ѷ	Ԃ�('�'|�+)<����g��Oz��5��e�j嵅�k�2U��� �_Ǳ*v
����^#f��H����hN��PC�#ƍȤ�X���@��vIp�$��u��ܧy]9		�"s�ZO,&7�RM&B��<w�OM�e�L���m��-C��4,��1��&\�k��]7$�g|T5~y���N�n�8妀�����Ж8��o~�dovv�­��㴋�K;p4���n[^F��%�:�=��H���yM�8����YZ�ڊ�˗�߲P���yyO*+%��)�Js�%��]��6_o�|����MOn��L�����t�ȁ�EQ�x��{�c���E'��'IJ����-�ٍc���5T!�=I�:�5��}�"E�밼�����~���u'�I���C8Qjvy%'�M�5�}%��|�z(�?ȫ1��p�mb��$�}D�$o���]�����Ę�q,�m*�Fŉ
���cIj9��s�j��Ir*��֛$�b���0!O�Q���G"Ӄk�6�4���<Q:�3�$`&;�I�4��7�ԥ<��#������)@��?yr;QZ^�oT�1���T�CY	9�,�"4q���Q�ר��SQ��??���*'�p��;�	b���SQ�}
�V���{�n����Z�[@�^���֋�,*:��=���/\��.�f=IM�J��{�>sÆ�qP��E^�J�[8���#���O#������D�Yq�p��~��q�6I8���ar!�SǪ�'qo�x�l&a��0d�xJ]��cy�jl,9�HA⺈dyW��r�ti`R�h7����������wČi�e�t�f�&�t@ZN��k�4�Xہ�1�H݁���X.�\u�RÚ��]�ݛ�bs�&��ƀ}�*��͏)QIޫ���i�Y
��O����V����@�&�A��9���4�c]d	߈M�$8���fh´D�-�5n��hK"�d0����>\O��m��Xl툺,�2]I�/�7���IB�%B=�z �$�p��0R�NI�+Կ��bh�i�ǇIR�h	���Ƚ�L5�ɫ"��Z��|^kf(�l���	������8��.ryq�/2��?���p�&�w�9� �R��`����.��*{��Y5�/XM�_��C�*��$����$�覠���  x���#f?YiI�Tkex��;�,�b����zJ�)�>�M��I�=�^c�C�hb#�ʂm"-1"k���G��ʊȫ��q��'~u.����ƍ7����]A�զ !$>�J�l����0�t��O�����~���Y��r�@>���Rjm����G�~mmm]-	o1l��E���."W���8c�MC�p�ed�w�o&6i�$O���o8<�m�!V�m��w���Ν��/$�?	NB�Zci�.ߣ�Y�r��J)QH�8Uň�#�A�5��|�z( %=�����r��N\mxKU,�y�=���v8I���V��R�'Rq�x��|�؈kp���4N׎�m��}#"�S%%<0���߲��Q������8��\!����h�V��m�6�#ݦI!~WK�WD���Mݴ��*��ȳHOs�$ʛ�3(���d�K�?L���Y����H؏�d%kV���>Í��>���|��7�I�B��űv���B6~��|[��q`&�*��6ܼu���\�	�9���<K)!�=�gy�v�&{�3g~D�撤t�q�7 ��G���~�&��NR� �%��.�b�A�&��ִ�m��`���C�Y&��:Aʈh���n{3`a fՖ���4rn����'&�>�i�"dnǥ:�;��v�Kޝ�'O>1P������{i�S����d��[�閍9���������̝�+T_Ϩ(װ�&*=-��=4"�!�T�2�:�T��$�aN�����٢G`#����<$��L�.��G�lB��-�]�T���*	��[;��!��W
��2:�pO��HC��!��p|�K�7NVEJi�����u�W��B?��FZ�D��L/���Px&D"Eo)vq3j@,7RU&�>�ΫKsa�yi��m���2?�a�Y�۞n�/�ޡ���f�ǩS�΄=w''']�^�;h!)��h�MF���_<~xc�u��ŻFQ�?~�tɑ�4�\Z�s�j8�.i��(�]��b�j1��*�Ӗ�-�b˦�>˛�Ns(�$��˽;�?C�5�R����Pd�(�겟�͗?�������o�$Y3׍���~g""=S�*�y@]z�c���Iv'X�onnn�Zk����dz��545�%$~��h��!�t��w&�<��u�Z�C����r�����]i��8��� �|���U���O�v,	)ֵ�]Mv����W�\A����ݮ��<�U5 �!�N�c�Iᶢ2��'��	�c�y,��wi��oh�N��#H��Y�� ��V�oDF����V���Z�y�Yic�����V9��D�ѣ��
v?���;�x}^���J>��6�|	���QU"���Y��?ۡ�Q��S���\���G�m? s*=��d)�;�w"��ݢ�Dcp�Ν�tL�3����T���#v����D�0���0o�-� G�����'~�V���x�('2[�qFF��pcC8p<+YW�e�];�|z�����b�赞�

��؁99&؄�܀���/���bAK̐5���[5��e2H�R�Ϟ�)44t�ə�>��k�= kk-ށ@�aR�e�h;v��g۪�o>|�P+�;X!����	�u-H�濔L+�*QhN}� �OL�c���X�ہ�T��{'�!��
Ę�a�0�#.��sU��:����2D"q2�.#+������*]�o��/B+#�dx<��g��OU��xO=�YN͌�E����	��

A���5�F��S�Q��������,*�����ۀD�>G��L�Sw�J?'yL��|\\\ijH,�A�&���"�~���v=�
��X^��b���O�\2���*��@���8JLL9#?J-ph��՘y	m���[մ�ZS��e����L YH|��cPx�!;Ā5��`̈́����>Fm~���\F��G7�� .j� ֓S��$!��� �����}��6�_5�EOe�`�pV��,�ʖ���i֘ �i�JI�9::�/*���֭���6�DG���w�h�� g�u�	Y��x���Ԑ�B~b�XzN|ej�Jr��{[GL��cW؋$5��cv�i��zN(LnI�sL��@��hP� d�WC�|���@�)��PU�[tOxS��,//�h��օ[�� 㝀,�_�u���.�c^�^π���J, �\�����+=}}��PUU7@����{�V�W�
��lSz��|�x��U7H��Ջ#����tedd�#h��(���Pl(���b ������R.�Ҩ �gQ:J@~�
�q���5+��R�zzּ��`T�?��Qw6�(�?=Kw�LN�`@�(۫I����Y�D�l�����BUj�/B@b#����u��s���UTz�.���S���T��>��}ܭ�����R�n`���Χ;�{�]|_J��8P��NV��������s�� ?��th7[�֜}��*P��?S����'�o�����ۋ����Q̪%�Z�J���d��'���0��֣��¨�{�|�pVN��= 3���p%p�,��?�G�c��~���y����������{  ��������Hi����b��X�@E�p�r�wՁ4O����������A����>y�ys|ǡ�WQX����� �Z�bd JK��B����kV��o�w�n�\���u-{��˸k%Ф::bڲ����_=G�����B3w_��+@�;#nݺ�`������y~��[���C�r�a��$�`���~mo5����C�� rZoo�9K����c��z�:r?77�Nk,�6X������W�Ԕ��G����$om��+A��y	�q�8�E ��a[.c��}�!�>H����D0�u��볏�vQ�0��ͯ���h�g�B�Ɠ�0�����v� ��SK�L�Y�G#�w���#diJ_��2��� P�`=V���Z7��E�oL�*!5A�s��X�/\k�G,i�K�R������	D�i4��Pz^eô,UI�U����@(E��a��)�[)���O� a�`-�B�>�-�T�B~R4��"y9	�f�)���i�	�O-9��W_9A��k-MM��8�Є���%�P�2 �ҽ�u�z��o3��VA9��1U [O]��f��E��ٛ�@��F4G;� U�yz����DϐG=�p��s�As�u�Z��*y@�21q�4�,���~>[:,A�jڥ����7/Zo�읉�73c�����k����E {r�$�h�VCړ��I�U�V�vj�kf`U�F�	�x��ъT�c�lA�1�n�3�o߾�I\Ɲ|?	`rz�8绮X�,��h"V�Ov�Ծ�-� �a���e�agg��Pe�֫t���u��9?�$���}�NG���Y@7
8��~��d���u=O�w������Oh��)v��I�?@�;W={13VG/q�*E����W('M>ɡ=@������g���u�"��;�5ѝ=P�����70f�����Ѫ���)�j�Wfǭ��/��I��-j-2Lu�L0��]�* ���	ľ�Ӄ�݀%ש�m�%(hh�*+��H7��k�ĭ�1�4/[V�!纈 ���6vv���X�?�a�Q��n�$�l@�t�իW)�5�;���n�-�!cO�� ����%	M�NB��z��m)��R��C�.���!��D��{)A�g£J� k?�������])�)���Ǖl�g��
���ů�aD�
2U��i���6�b��߮��҈�H�]�R��8Vڡ̬,���.0���7T�t���N҉��Df�H�����r����B�'�����';>������ۈ���xfcqq4�I���,P陃Ue�P`��%�cJP۵�%!R�O�4��H��ȀsF�t�Ò$k����K��~?��\�w���\%;:�C��}����2T�3��*v񈼭h9?�v8�k���sp}���~�uua;6zz�$h����M�%�{$N�DO��R�Lq��Z�v���i6S?B�lY{~��ǜ�ˏ]�x���WS��!�?��c ���G�0�1G�S_���p]�)�8V��O@�lml�� �\/�u(�~۰��o���
M���͸�Z���ΚY��YY
�������7ե����}����?���g�����|�F~*Oc�Z￀�.�,P�����EYr)VB��moVI;fm4�j��g���@��q����s_��'�˷�⦥�.0+.Z��}q ���F�(��2m�S�	���̈\ǃ���2��P�4/�;J]��A�#N5��fv��yg��?�Y+�(5��v�o>���@��m��x��-,�R�'�������{�� �DjZ۹ҫ-Ye2�dߏ�gdK����="d�x��I�u�,϶@����߲f9�_�ˡݽR��e��T��Kx"`��T��g>]����{�A�O�UkhxO�g�KOj��[f*&4M���4����NX!�QPX�<��PL)5�S�OjJ�y ��HNIq�f�#�EE� ����J�����6��r��y�왯o	U6�V�4,�z/�t@O!�P�0�PP�� ��=��F50�,�ݨm�\�%����B�	jCnQ��S;7nQ�>���|��������Pf�o����I�]��ѕi�(z��'f��i|���	�A�w�Ø��&����%b��^ ���j�ZBh��!��,��

@υ#��-�E��^�(�(CrRg��"�&�A�~���Ю���O�g�qu��m
 1l�E#o~D#)�Z&�{?�h��af�� c���r\�"� �7IVA�$+-�Ut �xy�^G���C�`�o�k���eW"�1?uP����w�T����ű�� ����|�f���*CD��]�a�/7��;�h��T@]*�;o|�o��s������#������k(}dI��`��052���c�%F�I(�ۓ�Q�k�$`�ÿdkV�6��m&$~�*dl�+wD�W�+�k�4U�������/. l><}�7�����Dy�#������)�й~��\�vє���"��h���pav���"�� ��k��^G @�`���~([3�<6����9�뮃��S9����Y��O�7B��t1U��N@��5�k�B�<(�`'  ���X�W'�]m=*��R�^�X)�f��5"��  �4��G1��ф���z��oP4��QZ��By'�Ҭr�l50�X�׀Ð����ue=q�"c�Ƃ����/�o���-WT����Iȟ?UiD�j�9�2�
J�r�@���4��������"��P�'ĮO���~��a��Q�
�1!����0���zP8h��(�a~�ڠ���=��D�O���\m���h+��.$��|��b�.v���В�SG6q���D��+��j�Y�����G���e� J�n�?�̆k^�z��)�j"�	�{�\��#U�5vQ��K�_ׯ��)��0O�Mg�Me�0�`�)7��d��{n�D�3�'aK@o�q�=*���̊Љ�0�b�!0��vG���w8D�����k�������&�^c�o:G����ˣy�90��Y���x�-�����	��=���̭��2�Z���*��[�5�/A�T�_o�=����^ ���O�G�W<sZ��o$����ǯ5U3!k�_4[��:9�(>�?ȍ攫^
��O����p�F ���fh�+��������W���^����k~��Ly$�n�\s` �@�=0��s��,�GGyG�)��mC�* �V�"�qB�Z��m���w��a1q0A�:�˨�uؖ��3�4 �/hU������ �r����8-��l�J!22^�4(Y�d+�M�^�SVHB�5*+��{UV��[F�����_�����r]]�㹟�����>���s�l⋞;\c,�ӛ}d���9��B�г�+f˃�r$�X���lV�~�����Q?YQ,�cҰ;ТQ*���R�Bv��/�yyy�'Q��0�m��O��.� �ߠ�j[�����~����1��T�*B�ё���Rav+	27���O���0�z�Y5S�}�1�L;^�3ˆ�)�B� w;���QU\�[Ā�\7��_��2����ō�T�O%� ��#��o3��ބ��ɾ���_� ��y�8�����a����DTV$E�Ë������О�I���nc������9]���F��%���9y����&��f�+�av{��������c̫�vW��t	9�E��'�~<�u�vt��x�<0D�����?�N���9�Q{)^�~��P|S���]>`$�I�ɹ�B��VQo���	���{1�/�k��3:::�/���}�����I l����j^-��`�4128�˟���`�k���@��bڹt]�O�����ׯ_�S�V5���	�CCC�	u;4QUIde��������d���zy
���p8�d�Y8El��
t��leuu3�}	���&obb"%%U\T$6]|�/**j��ډ2J����]W���~�)m�{K����p�J���Vښ��W�J�2w5���Z��Bwإ.Mܖ�i��O
��������VW�l���v�I�17][�n@F�2++��H<���N~d�]��K���c�q&>������:�iu����}��FI���eJ(��&U�k	wn�dV���x�1��n�U9%��T���c�(p/%Gd�(���	;�����wmy��e�L탛�h5��Tt^�re�⩍Ӗ7Y-��˖�l:�^���jְ�`ee%��2	�U]�y"��5{��u��J��ˑ�\���
循�*�P@J�ǥJ$b7!�?���?u>N���2<���L��sG�:�`ĺ�����E����p��)t�,e�X�H�2Z�R�T��|Te��TG����ġ��n���O��4�@a��C��P�Q�!��3�C1m�JDSS�H��*a�FZЫ��g�K�[s��4�F�RŴ勺��7�z���/�G��kH222z�4������kLyQ��(]�گ?-��KY��(���yTq���P��4o}���
�W���KPWv{�wKB9��3<�֩��|W
!q������@��}SS��
���!�f���69g�w�MHꡃ�����-,D������>ׄj6�����.�rN�y�Ǥm�>�:αa���go:a^T��A2����}�D�c
�q�����1q����C��)�Й��r%w�x�>��&�
� ykuyzE7m�@��=T��@�op����Ẩ��������9Q�}q
����l8g�t��o��$��l�����Ə�\3�&r'���ofȝ[Ӂ����𗖕���g%��,�ro�����T����'��JK�tʶ��b/�TPP`������P�p�x��d��hB��V��-;�*��uĸ���F>[�ƍ�s��z����J�?���r��>f�������7�A�nB��]����3P�������m~�
�K�ӗެ��`g�����oE�-�]���>o�\�7@Q���޹��41z���YT�Pq[|�+���w�Q˳1=Q����D���X����J\JN���W�ޮ|��,gD�?��(�ɲ��Nc�zո*dqn��X�N�h����ڧ!�Q��w����CօG??=@��S��%��>���-C�%Y��9Q�+|}L�Vm�x�8&��(la��D���q>�}��5��FȖ	��GM��}%�5����b���;����i=@��M\��Tmc#��t��ř4�^^����"U� pa���k{컬fq�&Ϋ�+=��8RL7+,�IF�{466R10�LLL4�%��(�L~���rW�4��0�+�nß��c�]��g�
��sW;,B��E�iM�}�:M��
h��}0����^�:��Ǐ�UVS{θ�T��)��w�������?J]��̉����e�D���l��ᆠ����iJJ�m�~��b�U͔��x��տ �N1^
�̲���`y�*ȡ*<���I�pZ؈���r/�����j;8���mA�ϕ���o����*���A�-�����qw��(Agno���x��VE���O����(��R1�u�gƣ���!�F�X�t���V� "�g*8ʼi�vNL'v� 5V˱����x��x7hG�x������@�eϠϹjjo_�/v���|�tj�:�����C�E1�`�^���(\7�}BJ�p�XS�������������o�/��0�2���������s555|���&f��V6pbҘ�w�v� ��@�vo	������?{�l+����E����ܐ;�'E0�y�/���{��#C�����7x�;���+�
(�H(�lg�%Х�S��u2
�d�����a�1.L)�w��j�%�U��M+q맷���WVVD�#�ܻ��|8(����A� ��N/���+R ��w�ې�n�&^��ݦϛoa~a���Ԇґtt�=<<�&&P�|����[ $ 2�^V��Q�at>�Q��N<H,�G��sssrr����/�;{�w��|��5vwo8O�h"���gA��~ӈ��^@e�`Q �/S/��UN�s��%�39 �nBn��J���;��:��)���3ww3C����8�9T͸��K��M�:�Z�ߚ��`t�]i�Hd`F-��]�cQWW7]k������x�J�����&Hy\$�=C�4����@��;T���ۑm�\P��`�kbW���7�7�4�x�.2��"	ג�=���S�����H鞞�����n��L��5�U`�a���d��m�S��o3�5��S��-#?�~�
�500��� (;�D�UM�/utv��O�� �FA��s뼽�t�ҡ�C�ng`` �Ծv�����M����Ɔ/���$)���O��]��k��nr��3��Ҋ��֒�Q��bW�p��5Y�^Y$��T�p�
y�n���;w�ܷ� �%�e��xҞl���:���E2F�w��qt����{�yB+	�ʊw[��/�?��,�0f�|E�3%�#� P�gϞ����E��1�3���|�ŉ�աx5������@�>���Z�#����u���wܤp�*ou"7�{�M��4���M�AJ��������Oʄ�л��#$��\y
-�z�����������W���վ����	��,���_
��I��ʁۥB���셬�^R��ɐ������Qo��8���1�nX�؍щ��͛�?�K�����:��W�Ǆ���nN����b6y%�5889����[�w�Đ�>zmbd4^}��Y
T�/_8ED� (N�%$$�#=}�4�r4pt,�ﴶ$�I29��n3�V%a[�E\��&���V��>Q�X�ӽ��`ue4a�;T�g���C� �_`�`�(j�Ns�Z��v$��&rbk���ٌ����' ,,-K��"'M�~+����{'����jd��ݏj�Y6�?�l���[��x"oh-���Aac��I  3��[0���C(�}�����|轠�`�S�Ay����2e�<~�]��{��FGW�RV!'�A�����!;�=�%�jW:k��8\ы�Y�񣚔@�@t�c���+�"�&b#�v9��pjh��f�o��^�w�$��������|cWX�5�Hl��9.�&���v����E�8߬+W���e��D�B�t�����!��3����}�gΏ�#��O�s��j$ߖ��o�D�-�\�	���ZX_OJM=|���w<Ӹ���o�=((�7XK��0��Jo��@�U8��P�;�#��ZD�u\�?��>�{l��Ī*^��6hN,���GM�+immMX�����7H(�HK�O������2������ �c/o����v{��������.M�Ak��5�xM����,���[�i��ɫ�iQhPVn�E�$Pr�M]�(p��p\�h��QPQ�L�6�iRS{��T�+))�a���8Y$�k,�\�ZK�g������;�*�Ht�qT��W7G���U�G��0�3E��^+P�����ؽ.d�YYT���(��w�MQ�F���*���������{���A9G�jNh(����zH���q��@�'�$�6�+��/v�" P�Zѕ��
�}�ɯ��<4�}����*��E�,ⴚv@�JJ� 
G��T�B���'�AA}3���G�s�E?i�uˊ,?pX��E:]�t8_t
�n�3�*��@Џ�͋&)l�V(���
12�"{�H]8��)�76�J��"!l��U4Bw8�y�t�#;�|PfGZ��-�z���E��"�DD6b(����A�8&�re4nn�)cV�@�Iw��H\L�pL���*�qd	H$��sS��6>�d�e"�	�)�e���!���P����8�@��
ٽh��~���P����%I����*��RQ�����E��Ӽ�Ꮤ&O���J�� �!:�Ō�t���%%�A0���l�G����ܔ��`�#,�et[����Kɓ��D������n��I$" Q��Ĩ蚛s;M{i��Y(�76��҂�C;�nP���Z��J9[�g�ys��$�&x�ʑ��E�C��gݗ�A=Z���7�)��co����8���84}���aI[�,��/�W-<V��^��n�y�51��΢���qT�/*�q�p�>e��ԕi�)4]|��&�^d}��b'V�f�-_VVW�PNM�fCk����n�)))�E�>����{���D��<y>�{J�o��8L��������Z�a��d������Y��#�[a�{�w�WƖ��^�D=��dٽ���g�pa}cjj�_]}�&֘746��Lc7N�sv����$����5�܅���W[O��R�T�KS?�+���&;on�;,=�^Yi�U��o��		��/��-�.W$�IQi��*�Rhu,U=J~�:�q�[CY�*]BSSs�c����ӭsK.�����V���7@�A=��rC2�"�C�j�А.�����c���Uv���*�!]�Ųq�iѫke�?A��[&����������θ�*�)��E�$����@���*�����Բ�΀c��u��$�i�D�Бz�jΊof���C�8��ބ&ˤ�x�Y�gXXX� �A2_���`��`�k�~����겎5dP�ۺX����w� w �Q}z3͕�&��z��2(\ˁ����o�$A�K8;;��a���N>�Q<?ڌ�F�ҿ81! `i�7���q#`+o�����.���'�Ք|�Z/ҸT���z˨H�_TTT �_�:YȈ� Y�񶎎�qqqw55}��;��:<�?��F��xd��c���a�N�-���5:hk3���}��sQkmm��\D�{�=�Up6�[������Q*0O��Yr-���KI �����g.����|�!�vzF::̀��p����Dc`�&7��z�L��@~�ZKq�� �������Z&� ������o@�K%��zO��v�D5v�(����g����ϓ��"�jI&V�k>XEM��>
��ؘ!T3-���B����o���`A��=D~-� ٙ`� ��s�� ����^�`QI���h៬�A�B2@\z}q#���At�8'��v[��I���w��J�f��,Lv3:::��0v6���x������E���6���$b��(р��ST�̈́�I����;�P]966Vܙk����P�.B+�u�Q�y�)�\���ML116.���s�x�8��6K��l%__%_�s��,iDԷ3)YY�H9w��]_?�Yo���W�Lj���)4�Q��%hC3��6.�H��b�� �M=�� �z�9As��+�m��jl��@nף�H���r38��6w,��G+��>��&5$��t���=n�_:Θ	P��F��>
�x�΋?��4解�a�"��螁ktt�[�:��X7T[>􂔨��v�JH�e�{�ZP2��V��*C�c��i�хJf�E8 J�M&����ʥ�/�} Pk�����ZZZ'��V�Gwm.h��%ݔ�i��@����P�������u��Q(�4o�#���Crj�?�4!����R�[����N�"�� �v�B�Eڊ�L��l�9(��Pȣ���\\����&0h<,!�r�l
�MT��8�7���ɀ��ז��W�ve\`W��4�{z}�z///�)��Ɖ!��h�A�"�9�epx�/�`�ʊ��Qa=@՟��}�~[�\�E�� !턷�W]N�`"tyk\h
ncf٘u��2����ũCp2��`�C$c�R�jp��8�%:��t��o	�a�]#�����.��������h���{hӾ�����xS10TU�?�Zp��Y�c��Y�r�X(f�[oq&(����x/AL+q���}��࡙��J��?,���M� LH	`r"	
R�č��5vo�v�ҙ34��08E������i�pь��_4.y���W�����1E>�*�Ϗ��OG0UVU�zqPm=MĶ����:	#4]__�мB.ٗ�l����0RH�Dq}kK� �! ��e�Ƽ-�����7tn2Q㍨�H�t!+��S(�FH��K�� a�U˷ۡ��{�dS�������a�� �����C�K({|ᆝZ�Я�$�ddd$�Ő���@�+q24>0�����|Ң�vU�����1-e*�F�{���A���&��B�8C�{Od��y�6�A�$k�ՕN� �w�����<6qS�=;�5�p�����������#�T
�ךlik�w�������#��d3���e������0b̾��@ƠG	=t�٧O���ǥq�S�	������� ��*��:r�9��kME�<8�
��	 p'(�!(nh�gv8u��~����V^��&B��^�s�NG��~�kJB���]�r����G��i�j&��;���w����L�����_r�(䏉���j�!�P텄j�¸qqK�O��6��g�F=��������넥]A0�`4��]:�t�x��IgǺA���z�����o�{�#�/pp�!$F��Y:%���V��dcamSu�� � Ը3��C"N3ҥ�����J�7G_A��U,�W�p�Ҁ�� h�t�G��j�M 2(!4V�{�=U�z%8Eꌻ����6�
k*�i���̸��ͣH�C�HZ�&g��K_b���l�TUU5]]'<����ߗg�
�����g�3e��=|SX�t.o:��32(�f��nQ=7T����		%��f�E�6���iP�}NK��yP�W���3�m��r�"h(���Ω�O������?A�CT�,?1\7@�q�	c1(W0x���cʢ���b���áw� "��٥Y��\��V�C(m� ����\�=zb��q��Q�/��ǃ�Dϳ���r�|qC�A��<�5�,�	x����?~t�E~l�GJ{�1���2��lmQ�r{��q�K
f&���@#֓];�最R<]Ũ2�oCn`H��yl�N<���E>V�V���ٞi#C�u�z��j/abbf�=Q-�0������lcG���6P0T����l]II�Ɔ��iW�	?����c��W�[A�11
:��=h~A@ݗഠ���]�yn���_���6����'̡b"x72�G8I�y��iq48]�����4:z�o���;�Z::�v��/,�]:��T�����ι��a���&m�3���J����9��.Bq�t@���|e�W�J���}"��<#>!6�;�AGb�1 *�ˑPgF��@y�:xSD�
��-yQ��`8��/#��h��lg�/o�Q`K��"�r����֮.(R�x:1�Ah 9Z���q>Q�B�m��> ]q��t�v<�������t���ߒ��M?Y����� V�����Bd�\Aq�GNJZ:�
q�!e�	Cؗ� �)(���^dm��z�s9}�yb�|��볝�vTN�w8�|�����'�R��d?�v��yL��(;�h0������
�1�r;Q�VG��V5���e�����`�F�2@6�����#uޔ��#P�28l �L&�\�v�]6GX7���:+?	�9�!>��I������QU`u�Hcvv6��{���Qȃ�Wv�3U�;��%���颭%������+�����UWG��	�6�o�����)�d/Zлv�?C�=��;bw����������X?uxS���+�|�SC�"�R��^\II	hN���{@�Q|a�؅A�I�����j�F������L=�S����}���L���1)���jW�.O�Hc|rZ�+lTz���ϲ�s���L)��V��b��:�m���2[dX=�%?�I�M���^j(�����kK7�5�9����][�1�G@��M�j��I���d�����.���Z�ۂ��:�U�:+++���$+�����7��B�=D��� j��\_T��qW�c��V��O����p��`1�b �a�I��^0�=��ȢP��[Ղ�&L�I0�5%^ǵ��7�~��%�!1An3R���`��vA	h'4�@�L��A�|PSOrC8�^��h��07���iu��`�`ܑ�LxAgҗѷ��J�`���ҁ��oϚe��"��E��%Z<z;�Su��<�0߷����9
&�m�=�S{Uh04(xW{W�-�k�U���v�CGS���E��~zn=˰w� Q�w}*��Q�������
��eTO"](X��@�`N���?��bN؞Y<��.3���٢w~t�q��7]����)�Y�h��l8_t�A��N�?[L����ڂɦ����K\�a �-���g�@�CR�[/|�1TC�3��bAae����ˊP;::�y �T��,�qu�&Y/���n�uyC�7V'c ���-^X ���ń�`�f��`3���3S�E$�X��j�c�z����e�j�۷"�T)�i���L�aN+�H���$���E��z�4�ʦ��9����mF���G��`!S�f�����Q܎��_���=di�}V"�P|��B����o1���	����`9W>�ss��1�]J
�c��dBL��x�O���t~���Ѝ�3���c�8lQ1cj~�Qzd$nL/�$DBJ����'�@oQgΞ@z����:�&��_hh[@$:�s#�v��?��/���n�-҄a���E�(y`�kQ��L\`T���6�/�:R�ܘr�����F�8n�QH�'bޭwn�A�6���7�����	��y����)�蛚r>��!<Su��uZ��@����B�JCK��ލ�����)���1aD���7�`��"�G f����Y�}�̊i��VV����`?�8^q�hw4 �Gc��}bh+=�����Ӿg��7�@9ޖ���-,("�8��-��
*?7����`s��MF��Aa�u�bkӑ�8�r3�Ss��(~ m{{A@�ʔ0�+�FX��sp��J�s]����q[b6���*�p
ӣ�%oB�N�#�>e�u�����Mq
1hԱH����3vqG�������j>���~GE֦�4���+'�	SfNNzr;������B��ނUP�����
�|!	� %������c�� Z�P�����C+Js�����"���-��in�'�m ��뾈�^�i,�7�&�B�6�މ�|��b����n�l7$f�O�	L�
4lpp0A�����^�8��	y���G�4�LD�3�)��Dm�#������C£84)ݍO�:�����_�gKF�Vzy���Z�ݽ2L���Dg�ـ$$�����S�����L9@}^,�>�}D�A
� {#��P��ܝe�%���z�IP�;%�uza.I#����,FA����[��$koF���1�K5(
4%'�����(�֢pp?�.i�o|�V$�UE�	HjR�_�p2��r`���]@�-�346��)�wuuE���䡥������XѴ_�5�ݼ~G�9x��|�|Ԓ�N��%s��|A(B��ZQP�&�]�+*
p��x��H�x�E#a ��(񥗠�A��̘A�.� ����h_ƴ=�SOwC���#Z�0��B�!��V�-��ZC"*��^�03`^x���޻��{_�sy��sg��6���PЮ�**��=F�����<$1�@x����&g�R�����D��A�:땶�w�G��X���p�&�̰�8R^3҈3�AAڶ���&=��������Tl�md ��9��NdOLL�n��7�Uc/Csä?]�x�B�-�\2?�G/ds�r���Ɣ����]��&$�/ɛ赌���������j�?4�>c�!�R
 ���b����:��ZrӁ��-�~J���U`ܝx�Yh���=_�T&�]�mA�>������$ㄟ*�UȰ���dn�"��Lp@��i��--KC�7o�D/>�&�������;�������S��cbb�^�����(��			K=O�E8�ߞ�V�*#����;�V^��GS:�K�-��-YU�]���]7�N��|{}���QVzU�#�~8~��D�2f���#�q���<Ӯ�/:���VKb�]�wN��J#O^��9�R��(u�)���8�f�j���d��1k�������&IO\��+HxC1X���|�lZ^�×U� O����YJ�V��~%!f����!s����u�?>nxv9R�wJ��<5$4�a�B�HFr�q"�㈗_��'͹�����<�#,l�ů_F��󧂌���J�_^�����mV�^�����)l7��Y��	�:%����2��#��;�Q,-��AC}}�9E���R���s�D���(:�����F����������. �X�y;;�.��E�(��� &�����9����� 8E���0+����[�>���hh4��}Tk���C�!,��9sm���T&1���<��I�}����+`��>'\�!���9���w�X��X$�e�������2oE0 &��e+(;���8G�=��P�F�al�ii�
���Y�ZM˙�9��Q�G�����Ճ�SZ?�C����w+++���#|]YYId����Pv>��R:��\"�� cmGG���̔��_500�Vp!nnn�� ����o�d6�p���b@�<���>��k-	b'"���*Vy�s����&�r�h���ݻZ��-�RS͕�냥ġ�E��K���e=-�$<����J:ndd}��r.!_\�ܐ�f$<��(uV[����<�r���b����~N�mX�	�?������/±��ۥ�����t�w�@U� V>�~R{���{��ͳy��0�R�`Y�7����[>��Z�E����r��
'�ko����,������Þ�4�,**��"L���3_��냙�<�4f��`�e萷8:�þ|�^�L{���p���p{�T�պf?�����c0��g�.������f�ıCE�o�n���T���fA�<�^��$K,�'���|^[�3�� j�`�[gfR��
D�WF����w��
���=�,y�����]���(aSuk��A�0����B��������8���5��H�����}2��q�Q�⁁���X(�R�F3�����H��066V`�J�ipSc�>�H�mu,B�������l�Ν;<�����onEɃ��x����ZJ��T����zz�.(f�j�-_e|���(�$o��ڍ(?Q�jik���K۪[I�����h&$�����`b�0��>�ty�|g��٥���7��N�WC�A���::�~85�iMi1�)�3=���X��r��X�����Ăg�I�=�{�;V<��c"���xx��3Z���Y��\�P}##�}�ϒ�k�8���LcŬPeUKh%Ði{[ٜM���X�n�3G`Q
�����_�lJ'Q�����|��.W����Y��b\F���b,��=eF&&�S��7i����V|,GXQ<�g���jJ'��gS���/�cYH���l��'���se8��
�	M��Lz"�;t*͆h�1M,.�rHH�~l'���{�?��!���ĳdگ�����x���KJ����#ƬY;f9B�4�/�7�hVh�"��?6�R���5�[���v�r�dJPv��]-��{����n�Y���Fo�f�O��E�[����
��χv�L��Q��v���6�y�7�j�R�9gBt���H����y�`��U�Mglk�>��턺Ї�7�� n]r>_��rHܢ�����j�E�;�}p��풀@\U�L���c�(7��;q��-3RlON"t�+�(2Kz+(3��sT?�߳9�B�q?��ˋ8W��i���tK❺�f�S6G��o�'�&Jy|����~RZ��1oIW��t\�}��ʧ���$�^���,$<[�l��*I(���+�1q��GM� �1�������
�Xa��={��+> @��̛��֋�x��xE�������QKX�f�5����8"3]9�)�7�5|�'���K�^����w�ry�����27�K�=ε�Z�h,3�z�K��#��ŧ�Y.5EMA�Cu�v��b�0�ЍL�ɯ]*�r#B�DU���$4��4v�x��rE]HO���Y��Ve��U˝����T�Occ�������P����d�Q�q�A�h醸Q�gƆ���#����2`-�B�����uu/�sV�a\�+�z^=%����~�\PŌ��n��%��O�J(3!������M�~`���m0���*-}v�ϝ�l�q<#�w~nn���xbe�p�imq�O��I3aAA�fK�������QQ%͗232(���C�1�HK{��ff����R��Y!�+�UB�B� �Z:b�j������}}}�P�f1�~3i@����y[;_&%-M�������sO����{���n#���
<?�A�C���&Y��h�14�F��$c�,~~���g�d�x�ӉB���^�G��ѽ���<�~�E'?�dd<����_�6�w�����3B�wI1</��-�o�$}����'�aY�����a� ��.�3"�j������!!\"�V�-3+r����dv� d�N����E:�cUmKƅ h\j����)]���А��DOu���XM>2M{�\qqq)�s���?_#gR0Q-�me�t�y>~������%�j�Qo���7�5M���O��0d��� �ߖW{-��Op�N�0��HMMͱWic?�I7��Lח}�ʘ�(wn,���7l'�	}!Ng:�q5-9�� +o��e��_~����~��Pu}[[��I3�y�t�X�(� ��|E+��e#��-H��2�q��!!3a:��`_�J������ᣚ�������ZFj211Es˝;
E�wY��ExJHT�R�Z�H|�Qgć$]=��k����3t��O��J�s/CU�c�>|+[����d�b���0R))o����y]���̓` 𡤤��I~�y�{QЛ=�b<��l7�`�끽�j��8�sxCo���;���W�����*��c?�0|?lÚ��-�ܪ�lho��;� Kl�c6��V��o��_�43��:��
���ǧ�'��K��	���{/ji��T���MN�n�z\}О�A����v���%z���=���1�%?ٝl$.����%�-�$%�ؒ�\Z�tc��=�ٌWIJK+^ĺ<�iɰ������^ ����=)�C��SU��!�#�~' "�Bt�14wt�U�=��{��=܊����E��b,_mQz���x[=�,*���'�5��5�헬S��gz�k��\��Z�O�o*��L����(�1>Cup�	�Z��su�2��*jj�Y�.��l���c^?��~�.VGS���I�s��]S:$D���1�P��{��q��o�C��c9�E�"TTU�u����$j� Ny��O�R*���c���bUkfr2���LHUQ���Y�-������X�� �ђ�6�h�,ls[9�X
uuu���.�v5]Y-p[�<ǋ#Ɛ����PQV�[��a��ߗ��i��6WW:p� !�&p��򰔙J�D��7�A`s�92�XA���ܯ� Ì�bqw��>����FNN>Z�:��s-�eb�y���WC�z�y�n&�
!ޖ��2��G|�5��F���R�&� ۗ�B��AvQ�6�h5�<z�訷8�a�A��1av���v����(��N���u��0�[�W�[��:��G\������=T��X����3g`b/@w BS�a	�G�={�bgɑ���N\�^4����qk��F9j�2vG��lI/�:�ى���3� Rd��樨�7�;�����-����n �PU����Y�9��D�7�
S���g?��1��wR�  ���|�I�,��]?G�'�{̾�O�����W�%*���s�/~�˦w�м�̃3��Z��kM��~|$l0�k�n͐����	���j�1�.]�,3S	�`=::����Kz;6!A:|��y.�ı��+�a62k��H�],&-�+�����D�6���q���>����w|��ʲM��SO��W%4f;��S&$�d�L8�����d}�`|�yv~�n��E�z���5�|+^ �g}6�:�G�
���=�sUG�4�V����qT�dFr��y`� �qxlZ��y\��RA��u�1S�6G�Ջr�����i�ή�WՂ��9��'��7_L�B֗\	����m\��􌌐�i�仯*�02*�����#W'59
�R Rï��%�pB�/��Ƹ}�0s�on�6\5�>d&R!F&��Hl�]�/鞃Zos�x�u!ܸ�o�?��x�Z��̥���ӳ�C�p�L��m�5�+�SDY�F�%�V�nt�^\�&�7��*�S����It�� ��3l����0�7�yp0u�ǏPF+�uD�R�S���6�ӻ��_�g9�](E"�� N���K�(�QW����J���<oE������
Ik���CGSf
V����P�ƶ���w������q�y�����*~���J��kkyH���\�f�f�<X���p2|ߵr�V��×��4t|����6@O��B.�`�=�'�؆A#��BTM�	vԱ�{h�|�^t���Y!#C�!@HPٷ؛���>��>���Y�Uy`ֶ����R�p�\8W �dӊ�/.�}O����1�w��u��A��ǽ(�Ӻ�~ԡLZ���`w�~�|�7�G�$P��pݙ.\��v�Ú���� z�6@���?;��-��(�� ��*?���Y��l�8]p[H���P^^~�مG�� R�����'����Qt:==J���@�wɨ�؊��賎?hʁ�>�wH��7��ihQ��`��U b���7N��I.��
�
��x���z1����1冚BIӱ�b�L9>>Pﶬ�/		IC}�;�Z�C.��]P;���'�[|����?�Pt���6w�^h�7Y��4��J��@aP?iE�42���f������94�����"C$s̫����5�P�=��õ�T^e�c�6�s�IBd���:멃H�(��ݶ��\m�#,Ec[��f��|;">�f��haUO��<e:ؤ�A��n�٭��D�����jV��<ƹ�p~Tj�oI>���d#�xЇA[`/T� �vTS ͜>\=un��=�{e�L��n�}�ؿ��fd,�?���^�% �t���t����R��>�@��Zu��a�=�>�||��~�~ݹ%�Q=�������kk �ޞq����G��\� ]4Jq���>~�f� m����1�e>q���4.���$�%A�/;���-�(9�+Y"�F���Wv��ǿ����T��T�v���'��!��Q����ʨ=��EU��a:��aYg�)l�� |A��~�晓�c��SUEE*��P�hn�#%m�_��+�H�`"��ӬPĽjW�)��݃q����iA�x�%JF�g�
?16.�z�
�W*��_`AD�97�f�fte�5��nq+��4��>��{־8Ϊ�cs��;x� �(a�*+��LC�����(��L�Mx(CCG�05�Ǯkl�w�p^+s�� b��ydhbb �|iee%j798D4u���<N�\���ڔ�Z�^N	g	"y��2��V�$�8:2���/G�;\?�r������䍐���J]�\��JKPDS�=H���ttb�����+����A���H��V�RQ��V��32x�ϷD)��i�X\��������	���t��:���q����4�,33�7#9��F�j��>B�e�g�&��[lj�3?77��xϾ�扣,�_��4X���

D�+4�j�IH�h�#Ӳk�;Ah�!���e}PD4��
'�����y�"�GD$��K�^�bOG��J�����%���9p|�8Ey�4|]�j�c����b���[3,��K���z�������ߔ��M�{�����3����~�)��gc��隙��C��n����-� ;��:�;_��t�{�'���X����Yɶ��|�Mgg�ys�8EH=kh%N&��>��]��Z�$OG��ȧo߾��6-p�)����哖�� F����~Ձ���F��x����,������}u�6����ҫL�r���@`��0񸆍���K@�����v�2�r
`��ǈKHX�-���uu!������Y��<�@Nb���I�.y�ß4���1I��¡q8�ؔ���@ZP#f�t��d�ț����T*F�W��~ffƈ�ɪ�����R��"�'��E�I0KKY�C`�94��3�OA#
�ң
<T_z����F󬭭G���FFF�4������ai�gb] [?����ly���8���|���D��b�n����\�ڐ,�a�����{6��WU�&>F6�QlƧ�A��Z�S����J�rq�IF`i��h���������}�ͩ �vA��A3 h419`YX���Ң�x�%i�ezJ�Y{ُ�Gv��u�u��q���4�}�MMM��u״C?}'jp�E���68m�LzON�OH���F VUU���N����r�΅WO�d\h����$.���\12<&�L2�|�x��9�ү��ik�
iȻ�R��������~��O�������8��k���ݸ:l�fAf�V��@w<M#�ZF���$$ܰ���MM�Zu��6F��Wd�Ӓ�z��LmN�������l�hs�Y�ǫ�LO����ұ����]��c�+W��ɷ��%�=����E�:,�,V���?1��n�UoH���y�з8����O�������R0k%!!qe�����A�ḻl`@���
b$rҡ�IG��bvu\TT��~�/uuu����ڻ'��h0!�~��aJ/`r�Xz?u�fJi��F�it�̇���`��z��z�����z���Y+�q'�f����$]@�(J��V����@{�������S��[}Ǵ�֦˲9M�ą������h���M�:##C��Q�8D�g�v!c4�b��(��S��������'�Y�W�G�L4kj:禧�)s���p�l?��gI�'c /����Bh��lR�D�� >���*jjBI}>�Ze��,r�[3@f��A^�L	����]hf.q�{����걖#�6L6��LY}�|�PW��.rB�k�-	r�\Xe�~�嘀S�)�0E� k����-ӳ�����1ܸ��22ζg���t0���"V�㰇����'O� �&�Wy���nl8�L�>=p���ňµ�BE4� ~�H�ݭ������Ϛ�v&��m��}���N� �AE����3�>}cy��.��W n���r�/G�p��s������i�N���7^o��E0Q��M--w��+��$��}U1��Ū<�姃��7(�(nj�W�����h_���-	�~�*��lh��,����� Ɂh\��x���3QM�CKg@�31.��lL�v��Ӥk��NG�>1&%����>_i(�R0��D����c�l��E�S�%me&�㝌�{Xb��u
� '���ƙ/�7iL,�&�ھ���˅�m�s��M�)���9Ki�ugc�˛��I��v���O�#<����MXA�B���8�c`v��Z�2Ѓ�͏������ݛ�ݩ��Ȟښ��q�r��呋���]	_���X��?�/k���)3��(��:������K��(�W�]޴Z�=�š����/*��%~���4:ON�}5�:G��{�W=x��-��t���Js��R1E�bb�kIN��Ϊ��p��{��R��+���xn����t7+��)��:�9B��C�iA�ZN��Iթ��̙��#C�R�y�������ЩE`�ȍ�±�b���u��/|��e���o�W�Z�C)�;X0�J_�  5�� �Y`�~�3$4Tz������h��&K �x�of�UV�L;s�% 5r]�}hd��B=�]�n�"b��ě����^�2{\>XO�/�p�/?������U����m���LV�] MEG�7XfZ]$\i{h�'|~qq1��V�H\2k:;��*�R�E*��C����ݬ�L����$	�x���_I��$VT����Sʠ.�}��E׾�6�����=ˤ�b�D�`�=�5|/�+���1�L�I�[y��/��~��(9qqq�>��aVIN����q��gϞͭn��t-�8/9~��)�[X�_{?�;)��`�A���­@&R��7G���]D~�P1��d��c���j��xᝐ�d*4�3DQ�FCJ�y�H�Y�n��K���hB�'�Y�iB��V��Y�J��.=��ο�:�9���^��Z�Y���=��ֳ�=��{�+�ӢEV����v���5h�::o";���^->&�d N���(���i`9L��?$"�W1�궏a����e�p�2����cv���N�����A�d����eG sl۶m<�yB�m$%�RF�1~~���N��iݘ��^�N���6�6�����Qm�~� 3"U+KK}��Cɜ^�|�wl�2-���
��n�_sm5�+R}~?ȭ]a;M���խjo���fXW��D[A!�� L^����✚o��C��1�Twg�h)��F���x�cn�ea3��V�ͫ�@�VS�=W�1[�6�(%Zn"V_V/�K�򼛛>T�ϕO��+v��!������י�������Q]�n�|�6H�Fz������|R2�x���2�v�{&����ì��/[��˫ԥ�ye�W�F����Tl����/_�/fa9�A��ݗu��X�=���@�� /�`|L䤕+Vt�F�}�m2[t����П�����!Oӷ�^��T��[�04���-U d'�t��C]�Yx���tR��f�J�)YPc5��@rr �̲]k��������R�ng��{�3г���H���]g%+���S�{�u�j���˭k��]]���
�9h���Z��~�E����P��~����$~���w^$RW[��������Bo�Ϗ��Mǖ�^2[��D�����?��u(�ſ��233���}��-fƓg��O�ך��>�����k�j�|�{��}zTz� �s5�U��?,����W��N���ލo���{{V-	R�q,Z1��P�DD1��B�T�#��܍Lc��:���+<�r~Oˏ������'O8�
p�y�n�֛fK����Ր>ׂ饾}T~�< h�@���C�� }3O�)z&�q��А���t�2H��7c�x���~��x%~�b����YR2��G�o՗I�F�˺�B��S^��`W��y��y���䏐�t�SP55�L�v�.�1~�-2 ����5�e9�YR��J�*�|G��l�6�Ns@MX����Ǫ�Ĭ�J����t������t�LR}�uѳ[�����,���l�	��@1ǽ����J�>FEw%V>���GZz:��C�E��8 ~�-�4褗����ֶR�_��nT��h���UE w���]��C?�!v>�n�d�C�k����z��s[��1Qo�<�5��_�	(*.����1V�t���k��FD�����O%j�/�@�K4f|||T
A���6��/�Q�XQud�\������
���n����@��-�IH$�%8�!*�9�uq�?A�u��	4��ޅ�S�$C�.�_YI]��g��gQ�@�r��
�PV��{M5�Q0�1��!I7�NI�RɃ�6�<�x��Zvvv�/���}�C�����QTTԣӑ������^/�7V���T��*J�ض�O|f#b�Zy�X���Ǡ��l�-�uu�ϕ� U��1����lr|�%ϽG��*9�����p/��}x�T�����>���Xy�&�h���l]Pv�\��#/^SZ�@Y�~�+d���t��0ק�Ŭ�[�8B��f͚5�����1�9�w~������Į��a`�i�*�3>%*3��~��Ԃ��4��*�"�MM�C��#TK�S�k�轭n�����\��U��J�.�jP,�����h�։V�ǿW�k����sr������f�̋-^[�>8%���f���D�V���!��_�O+**Z�b1����>�Q��_����g���v�C�~CƊN�_!Xn�����Y��uTħ�R��6�{��,�11뇃< Ӈ�QBq�q�{������X�<=#A��錭��!��#6�t����]>Y�4���W8Q�^	Y�E7���}���h��4L�P5�O�$�Ƞ:�9G��h唋�%nnn0�D"q�3�a��q�l��~�ePYW�L�ʚZ��ѥ?'��Ǎ�	(��z�<���q��b��:!��W���s�b��~�&7-��OnߌMi,פ����p��aze�U�.��¡L�	M#��F����c\��3��4X̽�Ƶ�.����V��K_��ж��w��&��{Oʏ�ܸq�WH�`ҟBϏ��|�����/���R�Fs�)�����r�	k��N�x�.�ĖKL "�F..��6q:,��z8��v:�Q��j$u��W^VG���t�D�}}^���܉k "��j7�?���ac�n~kz$�Y a\��Ũ�N��M8���%}�"�<�Sh��{�)m=@�κ��)��ҥ�k<�C�^�*fG���jV�����-�9@�E����Hス���ǏAm����Pz���Jn���#A�۸iSJ��j�i�Mר�h�d��|���e333Ә)����l�t1wN�w"�a�b~�g�t��|����ml,���~�4�KxB�m�-�ߵ��$~���c?��������=��|T����J���b�}�>�C�9� YR�k�*H��
���g'#����աq�.$���W�x,�VRR2�i���]5���u�t"�ENm�V��4�����g��p�Ѧ�"���8�)Z�B��ӛ�>��?�.��f��:���:�O���)�Sh/���=�����|����1�
�A(Gs�����zgQ���^ul�,9�n�~�0�������B��Ç����l���4����*n1{��C w���g�
÷��]�v�*���*�~|�

"�km�N�u��=Ŝ��,t$*�������,s��kEa	��O�v�:+�$m��o�}���ѱ�{����;��]�Gw<W���C��mrIގ66��Y��=i��:�H0�P<:s��`��dS&��N��ڨ�?1q���;��4�B=[���˗c�8�0I�"���nڅdY��q����Έ'O6@�������]vko�e�R@�I���*(�7�Q\^o}&���.�����H�S�5��Y(�])�}5L�iP���]��#;�w�ccբ7�~�Dgg��M�D_�h����RHTsg@�|Z�WE	 �!�"P"��\�vM0*H����6�F�_�<�o$���E�P�qM,���
*��+����&)�+�W�Y��U�F.�l��P|���T�[�FG�!oٰ���*���XdMŁce�WXL�
��``FT�f����Z�%��X\Q�_�8�Y@�Dhҿ�;i�5�	����Í�w��RE}�$K�0���Ϸ��ٛ�::��>�YI%B|�=��ܶ��0��&�7S�C��Ϫ��D~Z��8�,~�,����ɡ��R�hNʽ�:Ff�s
E#1)��]NZ�fJ���f0-������Z�xr�ӧ
L^�C��qt\�s.$w���� s����,�p�m�{g>Pu��صV��eܒ����4%�q<�t���^��EU�gve�������l��-����q�YN||�5#��O�[[/�5��
����m�\3n��_Մ:
27�|�����H�6.V� ���Q��e��F�u���0`�6&����಍1I������j$R�=nq���nxt��Kv*�kjjR/t�6bvoF/}��B�x9""���/j���|���R�:@G|L�]T���V 4X���<�t��#E�OZ��}� [__��[�wS 1������Ȏ
H8�3�65���:uwPYt�����t�BtC��kb��3{$���b��W�f�s\�,���&'#�M?����h=��[r_gō��2=lܾ����ﴒΓyw�.7��x߳zs����<��O����ٹ��'�f���_k�2�z�ȓ���q_>�:}�כKm��ٍ�ο/�l+5K��� &M�A/�v�e��Z�}�B�!�~o��5�ͬ�=;���E�t	ޮ��6T�O6Bexb��8���WUt�W]�b�ϟ?��탿C3�&�!.�{r/�K7H�H6̻g�H��XTL��\�0�1�hYhX�lt՝���b0/��ab����mTӼNO$�6��;�o<lڴI�wɛ���֢>?��R�&�������g�����5݃#���~ű�zw��*憫Q�<�����U  ���M����7�GR��7䲠��5��+ ٸ���o�+V���%C~<���DhI۸b�`��4��ArG,���f?����e��A'.�uX�;�=S=�������~d�P81��60 �$��<^�a5W�<V�5wV�%���g�n����b�Թ�"��^���G%�:��vH�A��W�o�� �.4���͛��Մ"��+۶�7�jI�����s�>� ���녚�����$W�U0=��F������{��N7\�1KEo����Rv0�� 0�\��Ӫ*M%�Ƣ\Qā��y�~��'�7����B,����v.Xk����j���F+�$��4y���BM��C������hD}oT����Xxcd؜2������孅�����������d��u�'�0������w�SbEm6�#5Q�r��g$�\�$ �_��X(27��'�Ӷ�l��1)f�ak"�{� �[9Ւ(0	��&��-4���M�����8��$\�i!/�9��:8:��? -zخ����yy�����������{5�_�*Iz�4<5ԭi'�fҤ�zC� ̈́B� �s5�e��C�o�C&����?�oMp�/J��-�2�Yfә��y���u+�����ՎX4�E���k����u����q5�AېQ�ɬ���<��e�MB�x��5ˍ�L����QuJ+�����%�o�OV�r7�n�4_@hX{"+;��g.^^���{�J�宵����6��U�����o�h�;�p�%i�� |`��r���Lw�<!.Vko�ת|�l��7%���N\\�4S2����@ݠ�X�|��6 �<f�k��3�%=%l�NzOH�e̴���HMZ�M�7�d���o�k�:�y�ff��=�e[��M�M:%iL���'m����$3C!��j���ߔ�G��4/����LP*&��#[�L[�|�� �u�U�;��{	B�0U?�iQ!��o�%�v�!�I#���C��=��O1������z999d ��V#�:�>I4�s^�о#a��Gž�<�Q�jo�#�B�D���ߎC\�m�x-tE�����"�����F��l��5ݑa��9�sG�V!e���헃�
[!����'HȅN���H����&���ڮ�v���P��TI=W��ۜ����$0���2���O��O��	���Aw��Z��m��Wq��s�F����*�!
���OW)	9gut�NR)�N4�ƊŞ�DpHXX�]��B��,�Ѵ��g̢�R'�$z�]d�z��qZ7��ll��1�������6��_� �p;v������t�fټf���>� I�9� ��Zvc��NـK��m�cŤ���=B�V,��-�'����߿���F߿Q��p3z�����|�351�hDI���ېEYXXl�]�J>�
>H௩L޽Y,e�����o�����ϛ�jo� �>�^��F�m���ݖ���h1X�䇢��4���2.��yr�ѴHک�|!�V�K�EFFV��<�tjj����WΏ��UyB�m�v//��h�������{'�"?��^�fS&靘��h�u���8�X�����ޓ����P��b�E�	;�~��� ����t��
to}	B���ӏW������_e>��G���A|m?�;��al�R��OK^��#1�~A��e����4_�$�='AX`�K3�$x�b�\��#q��3��=t ��
�������$�
�&ל��;t6�x��$t�%��ˣ{�Sp�h���>���% �?(s-�ԽbJ�L��q6\
�[/���*���H���*�hs<w�T�2�ߦ���e�"�����h�֢
��Z߹������/�t#;�˙��9��!���4�c=���if��}���c=}}E!�Z� ZH��mn��!Q��[��OQU�3w>$.���2s��XrTV� ���zo$��p%Y w�@��� �:�����f��=1118�g���i�/�il�T����D�n-m �>�N9��X�B2��ja[��"L�����%�J���O��\�����D䱁'`��Ā���/�{�b��v(?A�N#=:��h�ק-����қ���~��A���r�g��2%o��ܹ}e���tw	@��$H��s):���X��N��HKKS�Xв"�Z���*��I΁YP){����c7�y�c��D�����pby�ZrM!��=��� ߈Y���+�����F��Yc������2����@��������6/^���[����0�����9]\\^ggo�k�4�	&PUU��B��\7>���H�e�O!?<`�z��P��@h8=�.�lQ_�eCI:   �>��3�?p�^��v���雒r�7�O����`}���#@��\~~�S;#��橲���=(�!��8��
�%�w���{���S���$�w���;��;� @��O �u���ޮ��E���%� ������w]�zn���$'��#�h�]�Ҕڜ~�w�~�.@R<9���#P�Ԡj 4�yidd�U����Ք��j`��>A��[��AF�#j�!��C8L���*p%栍�a����w]�	� $F7�E����<�����Z(�`�U�fA��I�cp	���g;`�ɗ9r�|D�_/]�͜���H��RQGJDM:p/7�E�L���ӎ�v���Q�Ǖ(#��_�^F��|4V���C��y~�GHL���������;��]�=:���� �ֲ`�J�t�و�q��iH�M͏0f��"�7��E@�i�����aB(ף[��F�ggg�NIiSw�H~D�@��#w���'~3KE�p���X��#*@TK!%�5���!�T^F_f@��@&������,�ѯś�?�#D
�Ի
�84n6�#�IW���yHYzTy�+��
�Κ 2ˀg�JJ����D��u���@���r��\cJ��=߅�|SLR6�K�::���k�M�2�3��m��Ex��,u>H��@����@ ����T+��E�(f��t�������@�0׀oxX]�[-�V}���
K�6 ��+Qso�����E�Y���������fS�����U
i D�p��I~l.P�>�:V��\����t�[G�#��lZ�.̈́8�>����F�H7�8�$%M� ^������q�v�q��֓t�*I��*�<#@֐������n�K���Hˍ^�O�k ��W�R�fl�X&:��'������ad�]Uѯ32��_P�L6�ŷ�VVň����V�֜P,�eKǥQ��P�
ڛ��kH�sD I)\ʗ�L� ���n���S��߹[��n ��y|p22Ǘ�ߺit�u�7%K&:��\E�[vVn��R� ^ �|��ƿ���C��==�WzE�W!넄�>��1�V:���p��U:e
��O�i$ҿ���Ħ�êw��}�l-T���1�5f�K
�N1��zR�u��$==-]��d@=2�XI�!<<�f�./C��!���q�\�&�i�l6�������5��7�t��������_U�������\� $�E�<�]���"�<������t�廬d!�B��Uϡ��=(_Ƀ��^�'B�)��ucTkƯ�zݿ�.Giv0�Y	�--��`��F<�u`@Ŏ��p�F��^��BAY/L�y5J�|��-�x@���۵(�itH�c��Y+DPd�`F��Q�����q$�ҽ�%�c�h�&77���l$�)3�@��<���mX�=�	��sXpɐ�(��q�&����ۣbmpl��Dt�LdY�4Ru������:��)H���B���$���S 3��_(��Ӄ@/���$�ƅ�}�������MdQ2uuu�zrss��W>UA��V��'��s��ZL��_�ta�#�𽍖"����� ӏ���;{���Т_Z�z����L�i��������z�p�D{�ʻ�A��*Fx�/i[:i@��PՋX@�ԺLaj�f�A���ڌM��5� y����kz��~1vv�҈�f�R9����Li���+}j{�zbں5d�U��U~� P*d��VB���<$S��sj�|���r?@3���^����Ѹ��*:�����oL�h4��Ż�v����s\[O�U�"�u/��mP����/?�[(�$Z�����mT}�&�`%�T��e%��k0��Ç/XX����./�<$��$�M�':�P�zMl.m�M�F�В]˦PP*�
!�|/6cK����9Y��Z���'�6�'
�H�Kx6�~�ƿ>B5V�
�,�S��N\��zz��b��S�NA��������m��R,dK��h݉�D����3�\'�*�̱�q�y�[�Ys1�Q�A�(��8�C�jM۶��`oOK�t�re���c�]=��/�ӈ��6����c���9[jB����������Q��Zooo��,� ���'���(�Y�N�\1�Q�>�}�a�aE����C�Pa`1����X�r@5����Pg����m�C�9|Q4
���NCCw��!p��O�|뺶��MuU����V��]s�E�B�օPf�����WiƝ*�p�9�P�c����Pۻw/���Θ�������:G'*�iR��' �_�H ��L=�y��ә~
���z�ȏG�c�˰���2Ʉ�X�����󮀇 Ę��y��5��=$$� �����d-5QT�t;d���64����/��W@EĬ�e�M�6�'��9D�� �4Z�ԛ>�Ґ��ⶒW� �9��}����T@O�}R�����҅[����PG�S�w5��:��
��@��yANW�(��sp2����_��Z�	���4��
Ҏ�԰���;��37o��տ|�r�$��iG�n>0�}/@��$q�3	����Y�b~��Ŵ@��.���s���(��z��2��(��םṞ즡O�t/;�z���ʌ��}��95ONN����%�g�i��xH���$��t�4�����F_w����+��ď�y���OG&u����{�v��#[lA�`��QH�NÝ*��a�vV%Kq�Y��i�S��Y0�����pat *�rDq�66*l!�?�so�
�E&*x��;��èbho33=�?M��VA��ϠSȼy�" N��::��$5�Ԏ�L��hAC!aax��������
-�))�z��������VQ' 2���3�)�.���n��}Tcע/�@U���)��"�>h��0��w�m��l��}l��'�X��U����DQ@׀�燺��~f�� ͷA|E��u^�Իz�\�A9�@{ie!���^�9g!�F��-���N��V���m�����Pe�/נ?�EݧŪ $�
�h��o��Ѧ	�}[[�6-GA1e�Ж�7`����%�y�oDA4�J�܏J~��֡r�w��`�eAw�n�U��c�aO7��<H3Rh+
���$:�y�R? &HۈŹ�[���%��o��������C��h�җ��1��#	&z��h=L$-=�D���h&���Uu���9�!��բ
| |BϢ����������	�DM$C��qdn �3�M������+ShfP9i(J�l)������:����V�� ����𑲵��E2��xI���"�%�=��=��
��h��F��NII� ?��R~d�ٷ��[�r�Κ-��o[A���wݻ6l|���F�'1 �C5Z�S�6���NJ(Ix���px��+�6 %��_�~@�D��\"*���p�P�#�DA�~��̙3q����� �$�����Bݺ��V���`K ��� v� 7!�@?��}��IE���9#}�w��&d��Dx���@�/�w�}Z}�s�4l��!g�d���
=�C����γ�o�:m=�w>��}���`] \Q�z�"�� �@��
)�x�PA��-.ix�[�e�7�vȂ��s�� �����f���W���D����^DU[2-Oח��P�N�u���ٰ53�Dr���9h��6�_oq�ҽ
�/��;��Яs!G0x���iՒ�o������8��Z`��|XG`�[��+���Y�*v�*Fw�
,���m+����vvB����y�o~��l���$Rds!���
zO[-��W���&%GC" �!W���0Lu�F@��UY@��G��s����RT݃� �A� `A+ kNHN����`5��C`F[:���蘪	���`zE}�2y�������ޤ�K��������ab�A�Z�]ꍾ:ea��;-+k�4
|�m]�ȥ/R\�jq�2d����U�o�
�,T�� �DD�w��Ǡ0)�l�i�s��R	aL��i �/GNf��Y���hi���M~ŕ�U]�#��s�=����^[����P})PG|||���е�%���4A���谿���A/L��ҧ{n��� [��V���V2�oiu`c�@�[�%L�DFtA��\ 3h��H����}�>���~������6�mk�~�<�=�P��}���y���>�6���V�E��[�[9^ۥ|�l��X�~��haa!:������`���v5�b���`�ԃ� �4_-4�2���YX��W�Ջ����b@�M��!��T0`h*�c����㗟�[O��� ��7\���y;1O���X��TU}CCïz��e7?"ɒ�6(	`A��]�/}�xA���p����t5�p�r�>{l2�EŅ���̒t��/��M�h5��m���[����
w��/<��%,��7ȩ��&���=�F�y��������!ˬ½rBd_؇{Va�u܅&�5���fw��3kW"+�|L�:Eu$�Θ�>�3?�Q�Og))Qѱ�~��������͔���O�d����*������M{W�reZX �Μ�9τ����#�y3��M�,�#ˬɜlҦա%����S�h5,�:K���%�����深s�2�3|�h�V����c�(X}����%[Q zG4|M:sz(�;#7���A�8�h�8�]��K���,)�%CP;�1_��F\�8�^�uN�i`U�����!�Jg�:�Ƒ,C$��c$��^Dr5F�
H�. �Ia ��Eǥu0L\g�5��L��%xg���Z�L�4\����wFNM7�z6����K �
��;ܕ w
8��Owb�]
������0�>l���3�[��F���̓r=p�r��I�Ϛe��^��;�L���⦻���`��܋{R=	5p�r?� �I`�6��|�@=xX�ql�z�l��5�����Hr�Sn��-f��'�?�`�Ӡ�r�jue��?���A�Mw����,YƦ������VC�m0�P��П��p���:xă��<�'��I-�V�E��`����$�Q5B̳��k�����5)\P@�z�Y(���@�M'(�{�a̐��&�P#;��@O5��5�.V�F��Ƚ;-Y2��!l�<o�� ���&``���P��}Lj�,6�G7��;��)�}����ܛ�]?�3� ~�0�S��A��NO2�f� ^�d	�Q��1��la܂��:5�Ђ�p�B�Q����Hg;X�#(�I�,�U^"�ryբE_ާ�~yY~������	a�ˍ�'D��ě���n�7���^��bG�����%�7�~1�f�}�x����{��4/�bhc�'�lw�x�����<6݉��>�0�U��Ln#�}м [�aඃ�+>b�k6�d�~�m��}��,X����]�E���Q�o�Q���|�:v�(�K=�gZS��x��Jg.���0�\.���a��;��<Rs�9�`s�	�+�0F�B�� ږ>��C�%����дݡ����]�G��ׁ���8���@��9�3q���v)�tȶ���������J		=0OP�X+ a��9}�h����A�L��=A���ى�<�Q챫e�d�Ŏ8�_Q�I�Q.VL���jN_�7�=��+0�1�1��0#r �y`%6;s���6�[���+�n(ja%�b���0� ��-Xo?PhK��3��XC��8���P."�c*��jw �|�qr0=g��<��D���9Z^�q�8�1�uI�  ɂ� M{� .��b\�(�ԖJl6���<L{=�E�� �3B̯8����A[ڠ���V�A�F�Pg���A�0�!Ѝ��y��`�o�F����EY@:�X<�A*���C��zй�GN�1ȡ��=��������64��M�]n�`����uє7�O���d0�1x<z�P�I!xyV��z��<+-���j��G���!~@n+�ۍ�J��7���6z� <&�=�=���[�<�#��t.m*hT\[�=�6Nw���2kAL(�H�2��[��f�"��K�{Xg��,��)�A+`�3�rK.�� 3L���<��1���$�G�5�&*����a�%
3ʑ0иBἇ�\�t�� ���'���=��@�w�F1�-��߽��y9D���}�fl�ϐ���V��F&�̂�l�R.�}������Л#O�4�ڽ��]柈��-ւ��h�y��	���롣7p��!x,�ėNK;���z���Ή�)����߀��7���o����d�|��,������o�����?Tyß�m�$��q�M7�����W�v�(���(��%�mp���Zv%����.����)��<����1�R�25.����w���x�,�[������w$�R��@X%�����~�O^��v�����*���_ծ�1���#��9���F���,�o��l,Y�x���nof�Ϳ��:���������՛y����d!p�la��"�LK�:�I��v�\SS3���o:{��#:�rqq�`�s��U��\����w�ȴ�`k��+&ѻd��;��`N���І���C��&�ᶌE�mĕ�\W^�m̑'z�Z,�;z����&����f�u�3�8^��4�V�naU7����Q�*e@�1�
/PAGq)�-�w;,Y΁D�p��Jg�]���HB�}��gqcK�NgN��2|;<��eǵi��8g���4���ma�mÿ�o����2$.'����G�a
�Іی?z�ؠ���NÌq��|u��_7 ����m�9���^���#�����q���pM�ΞH����t��vVc�@�hÝ"��m��w:��NK�Nk����V#MK�[�vǷ�:��9������fh�yP~��ݲ�8ۑ%|]�Sja�q��Ƴ������#}a�7�3��mE�V�ZZ$U⒣��n罠��Pb���P �X/���FÃ!G�}�AA�����xP�]�{0�A��G�8	�S�Ծݚ%w< ����H<��=��u�ʊ����ߒ%ȟ�ݲ7�r9��P9T��n��Oa�5�!�ȴ�
.��~\Hp+L�6�nq�G��6�U�� �5@�G#XA&��0"����x���&���cp,���~���ha��Ex� �p���J�����v`j>�
��aj��=(^D�8FG5A��q<m7�m� ���Q$��ë��r���fl�0ƅ ����	�@n�	�����6�{���XW��~8�͒e	Lc�6�9���K���/��w��1�P"���k`���Jc�KnN��cx:� � ��Q__o����]ϴ`��v���?Y�$���q`�3fc-���i`w <�a
{ (�<�Jm���A��_ ,���n�%�e�EϘ��Ā�� �g츶�І�ۂk�!.߇��6D����6"zH�*�6D�w��:=����:��6f�m��D�������w������^_?�Ӕ��ǂ�ҟ0+7箯��y��E��������(�F�1�^� 2; 2��d���5�hǨ��D,�n��q�ȭ���]n����[,YZ$G4a�J"��Vk�� 1�� (�bFM�F�:�?`Ѓ��..lv���`dn�Hel����Գs0�	J=y�/=��a=n�`(�l#N���"�K�vূ�ԭ��у�@����"賥����v=�6(�C����{9@�W��a<A�@�ژ>3�e��(k�G��|sB�������2�B��`S� (9C1�W��NDp5Fp��>�wb���gG]]]C`>�!�%���b�3�][oς�bzр��J�`��w�L����T�
q��U^�D���Qah+��]�U��GU��]L2@O���6;�:���M~�; ��,Y�f����<"��Wɵ�}455���ߴn�q�EG��)�X6fa������bbډ(?��e��چ��xR���� z)y�$P`���*������	j�A��Sy9 ��0����R�|����� �P����c��)*6"h`��I��bn5����*�
� #ڸŚ�q��gv���-���P�ȳX�j|�k[�� s=;���$�`y&�z:,f+���0��5g��C뮑n�����c����%����|J��Rn�W��S�qmm�Xk]��̞fB�ۉ�����؟����F���c8}���|�Q��׌'�e�u���E�r���i�K<�$�Ý"�l���g:��%䌗|��Sd���c���D7C"����_$t�2��z�J�?}dE>�������Є�O2�����2���_���+�ꔈu���?+<
V���4�㿎��u��(ϑ�2��&�F��n5ޚ(�}}�ʢ��ݷ���V���\�S�^�����	��U]e՛(&f�O�}~v�Nv�Ԕ�?v�:^`m��v;d�jSM��#K���G'&���KM�.}�Y�<6�wf=�;@��j3o��?�N2��W�B��蠣�YV����c���7�A������p72�ѡΧU�5P5�ᨤ�&Y�ώ�d�mQg'5��Cՠ�i$��rO��믧����u�	h�E�'��1t�4�fK�R�k�{�>��A{���n�߄PR��$���I�T�W_=/�g�q`�{w�E>�LmB�"Rܙ�?��dN��q�ĭ#S[&������yǑ���\{��ә�C1��_�Y��/̮��aN=���d���=,&�!�a��"$�
�VX�ߜ"ߟҠ�����0q��lE�������h���T
��B�"�������B��_83h�DPVN�?�<�I�[��ş���*9C��Tiq�*T�|�����R�
U�lg`x�ƈX���t�r����x���wP�T�7v��A�aC�c#"����j�_�:TX&��hμs�g�Sf��w@�X#Z�/��ԟ��Z�P�i�y*E�"��k���4L5B���Kz�%�uӷw�7��v�t�,s9��WLE�7)ͺyvq����J�.?=���oi�xs���_?prk��k|��G}��a�
/+�C�ŚV��IDC��wޢk�2��ag�{��?Q1ȑ�����ԩ���mV�Hځ����>:S���'JL���3p�}P�O�?��zvh��l��=��V�Q-([G�a�\�^-ꬦ���u\i�@���-q*�z�2�T�Z����n@S�M�ۂg3��-)uFa�I؍Q��#���@3�pJ՞ZjW�����d�ԭ,���(��4�"�.�(ƻG�Ѷ%��c���,�!�!�9u&k�d�S�'�*�2�R��s/���zn"����Zo�|�d�5;4f���"���db�fMigف��$ܧ���k�f��>�x�?-)����I�y)b�N^���ՠb�㿨��ء��rxF��}*P\�雓�*�^v
��k9CU�.ػ�.�k���1pC�\x��v�eӡ�R��88#$)G(,q�Z$�����z�V�7L(��.���6���&n4�n]3���'�숓9�5rr�oRs(v������X��@���8ůT�%��o&>�S�0��R;�z�!�1�t���ܤ�
U\�a�m'��IԎ8Ǘ�����bQ��L&:��L�RT��_��F^�"n��ݺ��{a����xn�Ȝ�_���V%�N���U(�Dq�հJ������B�k��$��fe$��3x�����cмǌD��m4��Rg��UrS洄s��W�x���]V�$�H��տ�,Խ��&;�j�L¤���J������I�(���g�m�#F�|*�)�)��"��t���T��x�֦u�J�12��<�A�]��<�ϣ`�ie�'��W!�Lt~X���r���[TZ�ckB�ǉ��q�8#��Ó��s��?Qct䘼���JgS4F�8��w��eD��ΉC?�[iB�[tU�M�&>��^�넦Nn�w�7ڀ�o.�k��{{L��I���Pqd*ى�E�HjV��	�7����K,���E�k	�yo�L�mr/�-���Z_�jo�1Ev4�}�3fI���o����s�د��l�zpb7HW��E���eP�+r��z�)Vገ,�/6W�-)�������ɚ��Yo�?��4����(d@o��|�J@,{uo�h)�9�2@Q����ws�M�L�f�(�i3Pg�ӵ?ko��8�5bQȋ���Ϧҕ�Yv�r��HRS���ki�(���g�a  }��Ώ'Y�ޟ�|�ڞ?Ш{��M��X�$����K�����JN,O0P�yK<fok���lG�w���IW7��LH2[�Br�>���0Է?���SY�9�Q�r�VO�,����Z����씬����Ĕ���觢��r�r<�<.>:��T?��\Ú��H�g��2�zL\�yp}_1s�����Dt�K��3 	!5Z<��x���ZO���&��;���ニ:�}+u����1�T�<���/)+f�!"ݯrЎ�>�^��!2+͓�w&N:~DQ��T��)C��k��ҝr��UU�	��`B�wF�C�7yh�H�;�F�+�)�(�q�u�^�Xj��=�휾�L�0�����=����j���I>�xd4�,�)�lL|1����e�^��ߓ(u�����t��?��o�u���4��` ��3�&��b':x���'n
)^J쬾�('+#�]#�iYߦ�\��2:�� B�iTc���Zs��
/E���lg10��})u�a`D�Z�L!�E�J�O�� ���P����J��r�0���%ny�a8]�r���������0L�.+}\��?�c`�a%f��C�F.u�^� G����1Rg��r0v5ҍ	8�D|J��.�� �e`@:S��O�_�`@���������J�q��h�d�.�t�F߁=��=#:���Ga�?Ƶ�s���e��M�bYL����0!�<�R����d ��5�����\�\]�0��)�i��:ԟ�V�Iz���x�*��j���l��	�b`#=:V����g=��j�b��Q���<�~|��{��7�mUթv~ף�2�Ա�r������dz����NM�d@u�����b�Pg���ݓ\nka̾R8ձ(C��<���{��fٷK��� %����bf����K]�t�����qR�S�t2�g ��n�?��w�T�&yA��'m���F�~.��?�Ni�I���K��u�{oˀ��5iyq3:S?fy*f Q�3��U�u��������P�;��ș��Q�nC�72�zs������ݮ�e7��? ��>`W�-i\��:����6���!�7�m�����M��%���5�����c���Z�z��Aׯ��0&W��{���mP�7��]Kŗ�r2 ��rq�q���ͺn6O�̿i���#���l"#�?�g]x�e?���j!���z�VMjV���}#ī�|�^���K*��dEi���_�>8��4��:��`|w���	�K;V怳����(�W1��Qj���´��L�x���G��1"U�7��:�WԽ���ok��NPn&Z&5k4�;&��F�,܆����ɖ�3����rnvS5"Z�A�{�S^�m8�"Gef���.֐NsW2�f���?O\��;�_�`����
��4���F�)�,j�T��ԯ�}�3��a���Ru]���:N}�,�J�0\R�O��8w����1VZZZ.lN5gS��9���Z�=5<�;����;�đ�߇����E����Fø�/������d������s�����[�7���
�%zm��9�F�nJJ���I��T�ʹ�H��{`v��ѽ�\�NB�%�)�rr>2\}(�ִj�&��r5z�յ*��n��E`�O�Z��5N����@���~��ި���D)�)��oY7�j��rF������]��l�xy~�&Y�u�۝�3[�.A�ya��z��B����;[��X5�,�LS5����%5v�j�j�7�[�S�Sv�~ qb���늶�0�=������-w?�}N�p�	��M���2#�w�{��Ӝ݇�� �vt��Q��u��6jd���.��5i��R�6=�
���WIA��K9�YVBd�[�G)�#�(�{9W�UdI��fxh����'�U@b'C(u�R�r��S��,»7x��ʐ'~9:�fg��;����y$����:�oW(�(���yv9���Җ�Gmn/����6jZfZ�����	`�^r�F���̰#�U��v>v����L��Tg��a�MJ��+����I�f!⪄������i�I��bW�7k�c`I�E�C+�<�8�N���c�0^�p$��Ҭ:Ĭa:K��+�O�*3��u�Tza�d�3���)���AS�ī���?�t;Įo��e ;����k���mrl7����AkS���9�_��=71�$�Zu��ඳxBgH�a�)�u��R5�v���U=��[�f�FzY�s39��D|�:�\������X�º�:����q3J��x
�c0WY[{{Zyf���@�.^�¾Q/�O~�JcnW�Y��V�}O火K-�g)���,פ|Y�m�h�s�.�I?��Ԟa����"�2���s��F��w/.)�I��[��C�����B����Yi�m�@0W4�جW�A&�jC���Z�4�v��Û�1�<�D�ב_܆�Lx��*���5q���q���W#8���>_��ܾ�f,�]��G�c<Xte�i���:���5��%o2�X3�%��i*N\�-�%	Qk��;��z%o⽞ +QwD��OΏ'���#��Cuݜ�,�ň��*�JM��iۤ2;nQ��ab'�����x��db��#�������0/I�y��j�X%��q ��˰����K=8����`ͱ�׶�Ę��O����)��P��R��{�N�4�� ۵�ô���i��
�FŞ���"+�<��ˠ�o�o�T;s�N��63L�����J�먓����������"ý ��#o��j2���|L�C��`oo_�' zb�|·���
eѠ(f��n*ԡL�g��e�~2�U|b粰ӗ�9�2���/۫���8'yʱ1��\�꥕��v-ɻC���3_�EY)f�e����=����=����/h���+�Z��b��V�S7���K�gE@�!�"R@A�a	�X�֕Z[AP�%3!��HXԊ�7������|g��=��˽7s��O:j@!WN ��rDb�c�����Ȧ�0G��FI�ٮ��뮁\XBWxu.�L��,ۄm�߅�X�y3��W����_i�׻��ٸ��Y��v+�i;k��gd$O}T%�Ti;�7���]0Wft�O��w�J�5�����ѿUv���S&�nI"ҽӼx;�\����?ȱ�5k�d���C69��cUz���)l��&�f˜���ܥ^غ�*�N[����F�3��v�O�a�V9n�y��y����)����'�ކ�o���](C���m��{Yk{�禗w=ݕ8��n.����-{y����լ�Q��Ӕ����9G�\ࡴR)��G:�t|����e�&D�|�ѝ�;�Q�����.��
�5�YmVP��#�aa��d�֩Y��OSo�5d;�;V)5�cteI�n%���K���낌��C6��{AD;��$#c�_�ƒ~54��m��D���F��Z{��`�*��ȥjiGlXM�*�U����b{�"��	��fs��%������������k�g�+f���K���/���^�j�ϩE����K��s!>�/�/�j݉���k��8^��z�,���]WIxs�:B�q���dt�ő��Oޥ����'�����uȚ7��"��7|�KA�B2Ȗ78Gܲq{�$1C�Į~��8���v�B�u$=�I�<Ų�Q�w�,���gB�6��d�w#��_���re��<H����Ir(Rv+�Nw]}�x
9K�8�N��kJ��e�X}�F�r���*��D�֥x�؇Dڞ*A��s[[��9b�ӹax�б]�B�6-�ZR(3�a%��Ʃ���*{���j���6<��sE�A#���Un7_�k�6�U،����M��y?���|7�WP/�%��j��YD�9�=e�*�ڛ��;�mT�R��&y��F!��\���=O�(��>��q� G1A����Lk�������ӻ�kB���GtVd�_ݖj�B<��IcӇ�<yED�|º���TU���: {0�+�Я*OJ=x�DS��q����,x�m1:���K�<��@�3�x��6m�
9�.M�:7%y��[��-|�z��F���wW�e���%��C�k�ۻ�a���Gy��5�?8�hp)�3W��	��˜�k$��y{�|l9?��=�5�E�!��-ݎ��̎j}��@?���6ͪ]�����y�b2��!x��+/�$E�O�2�z2|Gz���r����{`���<��_1z�nq�/�ڎ�zU��}��������$[�/���������ks��Y�l���L������Ym���ԛĎ��o/�\hd�in��l9������G!b�#����&oN+(�إ#� ���\G���S������)���&�X��6S�LO!�X]�\I�����Ǥ�fo����eP���Й׏��рt>K����r6��t�ذYr?v���NӘ�@�<!�
5�'��+���p�N��^/��C���䌽<��R4� ���/ׁ��Q_�fɪ;y�分V��'�0,�����cǸi�Z�e�q�R]-2m�:�V �7O^ƍ�������<�\��=�K'��6[�_����������L�`t����f0�C��R�j�d��&E��c�o�D./��"=�hl�J��}U��(}��q�X8�xOc���!ٞ�>!M�J�h�N�(0G(�,$�񡬐�J�Z׍C�z|�Lѓ1�� �AY(�I�H�u�,q֥���B�X���m�bR/6�a��hm�k?��C��k�e��������^�7<t[?��uHorU��G�2�(s3D �3�rnpb�q:8ٖ��~wl}����5�c�
�����@�"KQ��P%�/O~��$Q/�w��<�y��tvǂ�=P�1��7Rk����z��Ɍ�"���C�ߙ����c�L5����=��O�*��̸oxH)/�
E���q��<�;���A^wQ^V0g��R&��@s(:{20G�xj��o�����=��yn��"��jO�a-X}12Y��L�K�����	1���c�j0#<Ʀ�LD�Į&�_*Ě;�zll������=%��iMf�a����w�s�6q�.�\��ԟ'���efG�H_�H�㖢x;�ĵlJ����J녲QG���i�4o�y���5Vg���O!_�Q�3V��T{fx� ?�ß���5�P��o�E��U)����-w W1��J�ŲQs˗9�uTU&u��<�(��z�`���7l��O���d��Z�xb*۴�{�{�)\��)�'[;���:�aB�Ui>�t��;�m��T�Ho�@g����)��$�x��ґ�e�u�=�&�����s�';r��y�AD'`�<d���EJB�;f=�H(��b�����K�$�"��D����vN/��XY����׋��8��C�f�˽%�#'�5lҨ'�m<���l�o2.�`e)SX/��R|͏���x�;�"Tẋ���0�N���֭���:��zFq ��]G���������w�Z�Ok|��W���an71������o�{Ug��
�}9"���!%��c��y��MᎵ���}�<�̍��(�sk�/�iAyv�Z�u��G*I�d�	��r�8W�.Pg�6`s�'�����:E�k�-"�r�[ ���s�����X9�S�����8�=��@:]�'�ZI(.�Pj����~����GDѮ��䑢A�h��4������z���F_�~��g�dsE�0G0x^�s)\�4����E��ѝ�����Uy�<Kv���y�D̋x;�!7[�^P�#���	k�4�d}��[݋�0�W޴��v��l}�\y�!�zA��x2�6��ƺ��%v�Q:[�=~� ���j�����T��y��5��~S�X�#t�����Vm�����K�&����������j7hp�+n��g�<�@�&���C�o	"�a���9Q�*�&+��,��8)��~`_k_m�Ȱ�΢�S��+�J���3� 2��J�m���h�}K�b]�Se`#�����Y˵��[�y�����?I
�`x�d��SQ3N�F�A��|S����ى����m�Zz�'<���BT��9ۿ�kc��;�*K�F�H,6!���/���9("��21������
o��E�~�f[1i�En�����aCD�!A��B�P�(�QTooRD��lT�^�}�
�|y{t�)�^E��8ޗ�f�#3LsĎD�Q�ݎl=u�1�l�ma��0MvY�$2�h]�O��a���Ǻ;�W�#��/�P�%{�����f��D�o��t_ $E�ě��"�$�o�W����Z#wҬ� i[ɞ�[�C�F�bu!C�/� "/FV_�)���P�9���y�l#�6�B��]g�p)����C�Z�\I[*�Eb=��}�6G��D�#ߚe���w5>��"2]��;��8��n$mɍ�ȩ]��Y���`���Yj�k� �ʔ�m�-E��Z�E0�ғ"�=[�?t��NA������a��U鈺�l�t_��k%�X@4A������Q �B����y�֓�Eg�U��go�e�}��-�����`��t��(s6ID�PF�ې�<�E�Q% %oDJ�C�_��j��Wp_��@��4y!�I<�/�<�k�-8�ҟH�m��Qfs�^�lYD��7L��@��]���rY%p����M$���1�m�P���T�^FX/�2�E��K�*ԗ����G|��v���Ԋu΢6�R��D��v(���G��R��FR0�9�%f]��5�.���靹���e��C���O��
z�㤠l�x��Z�Q�Ke�AE
W᎑��+.#-r}�Ґs�{n��g�~��ђ���%㇯����ﹿ�\}h�w"�J��Պw�SG��������Ӹv/��j�<\��k�!1�='t�����2ǻx�<<���?��p�O�E���t�(��M��?�&��Y�MG��&ǎڎ�!&	������G��È�-+-�o��.�o��ָ�YYI�]�Y7R��MN�:�_�1�tD���I��<��l���7��z�U���r�i�#j�l�buQ��*a� lo�5r�iQ���:�`��*��2�ʾ{�f�_�M	�݉}�LZ9-�m_���F��W����#��r��~{�N?�5�>8H7�7W}N�u�ٲ����N��ŁX�j��E�����+���c�:���� ��w����<_X%�����/��X�������= �v����z�,�� ���-��EB�����b;�D<R�Q"����]���x�҆�MT8&dT����&w���J�����D� �pn����%
��1@GR޼\����hG.���V`o�8n7� 
��7@NK&�ũ�3C�;����A�]��\ތ��k#�6��p�C��)=�)���
;ĳ��@�b�b�J��]��x��w�t��O�#�b���h�*܃��0�a��M9���,��?���Oq��zѦh��zn6،W��G�D;u�'�X�v���唂zD>��?!��m<��ؾ�m�~�Gj�[��W�R_�<���$b��s �NdJm�s�����e�"�ђ�D�U����[�Y� 6d+��a?� 
9O)=���&�U˚�lݎ�uHhd�?���"��Ȓ��9~*�=�8�͑�&�����H	�ž�B�V�]��S���s�Q�[����2^�٣]�k�19}r�����:r(e�^�W3@��Yӌ�L��Gz���T7P���5x���[,�`U%��*�As�u.[�v�z�˗-��:�Z}*�$cq�i��o{����SK���T}�I�ۦ��C�T޸1�� D�l�U���n��*&�������S�ۢ*����7������h��W�����)���HJ��i�5
}pT-���e3ƶ��I6���kp��
�[���؍���JuTY�O���	�[�>^�n�@sZ�����?O9�$�]/cZ;b�<]h�l��!d4@��{�����2~چy��8�����nha��YI_�c���Rh)�|r��ܐ����#���R���$�G���`W�v�y��eH,��ڲe�u遃H���6�'�0���5�J��!�8C�.��
��lC�9�0�	�}-��d#�Eٚ
:�x��(�~���S�ҌH�^q��Ą���p��c�����@��*֢�_GM�6���K���W"M�B	_I�İ��
u����*4��
v���PPXg�H�L�j/#g�s�Z���wD��|}1�AK,F+�#�JjĢq�m��
�������m�OG �\��,��RЃ^
NƟfD�Wz��^x�z!�U��;���r~�=����t�qҎ\�������U���+m��v)RZ��f��@��_��L�.�[G�aǅ��8�E��xV�"�V��U�$�"ϼv���p��!�_�q��x'#��E����\f'�_y�Opp�v!Z�GF����\T��[��v��O�v,�M]��zq��7��]�S���x�o2��i5���~�]�v�,�q��=�\@���x��<_���N�A�����R����p߶Szj��U��]�\ND߻�O��˟�W$45�.\��]���~�Tg��$6��,'�G�I�r��L�c�ωA�9�:G�C� ���3M,�0ݩ5H�ޤ��U�w��uE��|��vz��P�<�o�c���Tl)�Q~�l���ކ{�K�P�A������̃G�v��U���Ux�i#�el�Y��RQ$�%n��x�3�<����Uu�Y���+\\��R�/�Q���@�K�{��zZA�o�ޮ��f��2 7�`T��U��0\;��
-$���TH���]0���4#��B���?� &Ըq��]Y� b�Ĉ=X@����{�
3�u��4<�5�d���U5��`O�F�,<,�kTCS2*�Yf��b{0&��M�^'��.�@dg�WŽ����I��u��3V���۪j���N%F6���iʟW&Y��#��ۛ���ɼ�G�%�$Fv/@��lG"����K�#�B�ݗX��&�n�\DT���|�^(���yQ�3��V3���PQu!x�?���f3�A�z�w�&Uڒf�aѣ�.�V����ƕ��r�{I�qj,��~(B���0�Ryܦ4!Ʃy=G"YUH�[uƉAo���*ũ�I<�T�_�rـ�[���]=�V��V�����#�Wo���ǽz,�+=y�]uI���4Y��ǹ��o�'�-�kqA�$S�s�u7���D��O�X�c�B���ϭs�ղ)M��~���QBl�OꟌE�fC���,�VzcF�^� T"��v 9G]�6�}@�gVD5��U�.�9}Ű�F�
Ծh.�;��r���u�8m(����z��Ge�|���\d�D��r�	gۣ6��Q�b���H�����"+k~_"�l��Ȗ�әTH�(�c]�������0���[�g�x`�k��)8\5��C�t��*����ߍZ���\T�N�#L��I�o"w 5��>�D��|mr�K�S�������-h"���(�>�i>�d1�!���]6r�+�
���c��l�J���t�B���OX%�!$k��s�?���=]v^��a�ݔ36���.tw� �DH�Q ��U����C uM1x&��
r�M�\K�yj��u�N�ٺ�*�HU�L����r�8Q���\���b�3�?�v]���2�^���Ħ֮�ф���I����ee��벳K�dP��B/�!?]��&o򅎒i1��!�":��-QfH�b�֘Dċ5��f�����ش���^�����k�"��3��T�d�����~��(�Niag��� ��V6F쪮<
o��ȡyaO��XD؀?�FfDv��SB}��nL��#���D�q>����Bn�l5e�¡�D�c�҈�0�Er� %�������+}���fL�[*ۦ�};�:1�EB{�#j�&��ʑv�w���g���x�׋rĭ6��]� ��uNG.Æ*}7A�����s��}�LX���$�£ŋ���}B+y�.-d��T~��F��:�e`;�mV-�a©�F�J$�[����uK����m'D�ݧ{�a̭ƥQ՛s�N;B�3��j����2>���1 �Ͻtq�|�X|w�㟛�xr�TY�������|%��P lC��.3)$����^��Nb~�<�=*id�i�nd��UeKx>ԹI�t�"ד�rh���M�Z�]U�����U0�p�/[U�a��~�*S�G��.A��.���K$�X�|gD����k�R�)�&O[|q�w�kb1�in�r<L&���8E��G4�VkJ�&�^c�����m#�2M�Ew
C�*��+ݕ\����D��]K榋$^-5M�1�=��#���a1Dҍo^�cX�-�Co�!j�s���规��Gx���lI����)k/S��� W��{�E�*��h��~Dlo:��(�"M��h�������
m�`�I��RE�b�UuP�o����0�i(6��#'��5d�I݀�s?��W{U� ,�VU�|@�*����+�]����S�,����r��\ :GŐ�x\�^C�$c��j����W*�6i4\��{�����|M~v�*�G6"�K��cYˤ�ċI~��k���rrE��)��i��|�ZB֘:#�"�H�zMӐd�=7]`�P��K���D3��SV���7�&��S6s�Z�KG��h+���|�w�����f)_�s������I�����&����<2����׺z����؁H�qC80;����rF��L(�݌�6��r�e��^�z>���w�J��9���
:��p���dFBt,d�1��1#��,��i�g��md=��n�.G�7�{*��_~n��ly��c�A�&��z�/z�q�ŉ���9C#��g8\�5m?^�Iq0JC:P�@�mg=�Ƞz�Y/�3(C���A���+S"Y(�%d,XT� ��@���m���@y�E�F@iTz-f��`P�l*�r,( ]`=���
f���[Y���_�px���۾��Ȗ���t�	�Y7�%p���_t|>ޡ�!q@b[ k6�E�i��}��X@�5yhdBgȊ��:�tt�����]��`lN���/�
$�@M��d���=���KGZ�[�tX*���~�ʑ2S멜��O"bA?1F��N0H�������L(�H`�,�L'�Y>�H�r��:z)��� ��9R�eS �2Ћ�P�N`�^�7�Z �Ӟ�`��Џ28��~�o����xM IsA�
���z@e�ס�^�@���FA�^���6J��X�!%���]����r[��7�!!$ƜaL6~n����4۱4�����.�jP�{u�w+L\���E�Xyy��Ɵ���WCUg�{%��Zx-�J+��ZBs�O8��.�i�����?�eLǧ%'�^��bT���1�y��mF�4���]pu���FX,�~d`[X��`�F�f�ʂ1�,�Øq��.�>�X�V�_�Lj��}irh��!��>9Q�S{D��1=&%)�,S:5�q�ʑ�	{�>��n�6 �,f�- +e�΂l��lBg���j�ME��/�ě� �8���H�T ��R0#)���p�Mt�Ft�7��m�IFtp�2�����8�-�����T|A��4ͽg|�e�:�B-�4����t<0��H��?���':V|kdv�?���J�t�q��`7c�:;듟���� �ۓF�s��a�ǣ�FR)���-�n��h22�ĸ��P�s�m;M������ �m|�E0'_u���;��\T<Lw�������`�DEL(��f^�c\m���+� ��Oǀ�Mz�Vu,C@�;O�p��M ���`r���
~+�$�-��Z:�Rn�k0��3:eB8P8w�NS�gƅs�н���J�]�LHt4I6.���ӝ�|���h(:��h-��e�J�ke�o�ŧ+��
ş��`�Q�vC��@rAрQ��5 ���v��g2�0�p�s�av*H���OK-���`�!��Kx�w_�孍��k8��-�5h�`�c����44�g$������-&3
�f ��e�{���k�����i3_f��з"�C�|8�����į4`+A��v,�8��3�b�q ��'�0Gf���eƁ�ǟ6�x�8��	ֶ`��_��-��>n_7j3t$ �m5F���r.���΂?~�5�j��O�r��q�QT�����Qmw��	& ����/��5�3!���#��	G�m��杦�F�ݗ@z��{��Go�K�L�H��K���ß�- I�	R�$cC^V�$Y���?rC������޽�d޸����po��?2�[����r����PK   ��dX��_8
  3
  /   images/57489f55-55cc-4ea4-8258-f1cf3d9c722d.png3
���PNG

   IHDR   d   .   �!�^   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  	�IDATx��\klW>3���?�vR�ql7M���aBih 	�F4��hS���H�

�U���u� ��[�(!IqS�R�j�4&�;i�:[�w׻���|wv���cg/�u�I��uw����{�w�4`H�b濙%�k
�ٟn�N�W�éR6���KCCC�v�����$I��$���|�aM�<p�@ʿ�Al@2vPq�	�L��᠎�jii���2ڲe�,��,��=�}��7�~�o�.>��~��Cs���\AY�)�1::J�XL�c+���b����0E�Q\n`6�?a�Z̜	[w�\��4�
�"���(JB��|>��}\��y���y�j�̝�h��t1 ��������X��rrr�6�������i��̏2�j����ee��UUUTQQ!���A�Xyyy
�(>ȧIp�bA� Q�������w�gQdvk޴��;�oN�G9��9c�ڲ��1��Ջ�x��^E�2�� vݫ���vH*�Y3J#
��Sv�y�F���|
!HT��By,�|�{�1J��i�D��O1ױuT�y|բ��j^ՈcwH�V���RJ��@.i'Iי ��L*H��ͤ�wyh��3�PN�������v�j�**b$}�O���#� 0ہ�����TZZJK�.�lc� �������137~��	�Ht٫ju��+�Q%���3�|��a[Hz�$������Vjnna�֭[iѢE��OD�@�c������������Gn�;�>�Z*�B�QP���u��r¯�����cتjz�p���OИ]�/3_3��_�����0��3�K7!ǝ�xvb4O`η�3��"��V|ְ�y1Q9n�O4M�.]ҷ
�"�"��0�M7� 1�a�$������h�8.o6j�0m�{�<y7P���'�lo&c��Y3���#�1����9,b �:Dzd���drG6� ��O7j��41NG"#�L��Z�4>:zs���H�̤�1�!e�?�>�|��b\�)��{|k����8v�#
`�:��ac.$a1�1Ě����2_$}�`��[�P
b��LwWf!�a	��T.m&� c�
��b��(�1TU�'��nJ#YɎ@" ����I�������@�������7m!�8�m�9XFB�|�]�{�r|����5 �h���T��)�!_���b!L��_YYI۶m�ˮ�>����0�}�k���N�ec>�l�J��'_M�ҫV]UN��������~����w���"d����.^�H�+J� 4���Lit��g�-[�M�����A!�����g�v�|����vwM�I�i��)~�9��(+$g]�k&��+W��,)�U!Z� �"����療��D6`%��� 񋵩��O~�܉?z��G���X ��$)\��˺�|�k �������^��h�����C�O0	h3�w�*w�o�N��p�7�Ap��W>L���p��OJ͗Y_t�|����Q޾ig��o�7=!����?�)z ���ڵ�x �or�Oix��a���YN'k�厰�dG؋��\�ѣGi͚5�v�Zۑ�b	�+ H�����-̳�=��)�03qc�AQT�V�Y# Az{{EZ�������S���&-A���I�:YǬa��|��i��	igS�l�1�Ng��|�t�YA,�Ę���Ux�՜G�W����kMY{� v��g?G��g��lG�$��q��MI&K����l�anX�g\%�*c>�\�<��,�F�)D9����R/��]���q�6� �q���"�W��3_���K��9tn��w�F����6�m�K�u-����`��XS�JЩ���1B�G��������n%w���HԈ����{TRT�R��DR�����yqu�0�G�%^�1k�9���+�]��z��8�̿zK,�~�oJ�EXz_گ���JJ�"�d��@�ŋu�m��wۘv�iqa }|q>�t�q?q��v?�_^�����>0Ԑb���Ⳑ�]�z5����e%Is QN2�3�ļ/Fr�S�_�i YEx�~���2��,c�,� �t�b�!�!������"�z��5Q"&Ǥ��b������ҵ@΀�,��&����s�GI�X�e�(��܈��+A��X�`d���&�dd�/�L{�rB��bx����DVbĳ�R��Ф��7���Q�$eOrр񢧵1,���/��%%%�����l�̉ �P��������K�:���6���Z@�c��.
��=Â��g���O/Y��������]�Q�E�\��46�]̇������6k0'Q�}
�Y�v�+W>��Y�h�U��7���\��� ^��z�ϝ:uj!��9s&�����d�?�`]�ḣ��k��(�ǌ�Qbd����-�Ik�S�l�C��%�KX���Й��%vO�g<���شc�aM�a�}�=�
�7    IEND�B`�PK   �dX�A�x�L  �M  /   images/6470d57f-e26a-480a-a2b1-cdb1a5d6cbca.png��c�.L�&|�m۶mϜ�m��m�6�ض}��ض���c���ɷ?:��tR����H%)X\X  � #-��4 @�!��u}�b�'`��]  X��3@�]Ӊ�[�q��rU�m��a�l���`�v�u15v4g��l�}͏ �Ɉ���ɹ�
�S_�.O��ZO�,�Z��N$%��U��)�/̟�z}�	 U��B�AKJS���5�6�z�O�lzS�5ٚ�=���\�:NrN��R^����VV$��eP�̵����샿��Oj��2d"�^4-��J��(<���LLL�����7/�����>��=[#��]
��;v�};���3nZ�z�?r��Z\,���V�����s:NET�n*~����U����W,X��B#�z����ͼ��+V���
����^ouM�<�h�����/�.���Mu���a
��G"�u[o�I~u�=yS�k]7ce8�|��)�q�xZ��{����-��<b�>a`���� 001e}}}-%g2��%+C�@��Qw�yq>����	�� *���͒Mk{�u6Z����ܕ���R�1��>�n͑�U�#�S��^�ԯk-��xs5Y3�38�7Lsj���\ߎҁ�u�Y�*��h�$�	�B �·I*��ky��]ڍ�_�r�YcMo��������k��]����n1|ب ɓ!��:�@]�7��9u�
�:7�s;
GQȥ�䌥 ��#�憙~`�� �(U�o)3�Q�*wN����:��Or}��քTc��_\@X�gT���{��:/3�ɍ�ID�H�~<_B�BŁ0�\���k��l#��,�k.�1���&C��� ��b���N�r��F���߬����8=s0n�+|�}v�ҫ�8�	�@�T)�ڰ����&ѱ�_N�K��yԚ�NPb*n/Wk����~�&s�7rFL:⦔�%C�n�T)��J 0��E��5'��jp�������;�:+�:oi'oO���At�j�>�P�1����mv�����Ei��(a2%�2�q���&�%2e�Rxu�������L����ۓ�V �Ra) ��-�^?�d@�dhPw�1(5�"����G�CA��=�G^F��Q�i�;�ϫ �Ɋ��u۶gw�<`��EƁ�\�-L��v��xH�
666���lmmv���#�ҵ��/�?]��GE?�{;:ޮڮԼa���1v�x_���g##�E�3u���3�d���3����S��NBa��;����U�X�3ge��n�p�7O��G��v4�XF�,C>�8�kJ�>��t��t�*����O�h�� �A�w8,��8N���}��g

<������ڮ�����Qp�B��ջJ:�6�D= \��S(hE��<����X���ҍ;���2(耞q�����z"+W6���Y.t�����7����W���#���WG���wM�Ht�[��4;�]��$V?�EM�%.5U�Oc�/�O��G�O���	ݫ��@KS��x�Br��k�M&H}U*56/Hg �I"*�i��-��j�0����& �d�B�f�ٝB��Z�����7��8�B��eI��LX�]�p�#G
��Hr�x|N���a���|�ɺ.���V�L�������8�ܙ,M �2��s�Ȉ��>�F"*��mW
}E0�0�3L�d����]����_���x���e��彲RTD*�-��ۯP���y�b�*zIn�Ar�-,*��A��T��*��軨����;���-�4�p�b	�TG#�;*�4h��q�%w��b�@IC�@ַ���F����� !}�׋��:������i�f�t:z ���p� 2��Y}o��v��{^���CO��*�s�Y<�S��;M�r���r"�˪_��R�����йi50�h&�^ɥ��*�� ����̫0q����1���QYB�����?�ؿ��F�����(I��M�s�"z���TF��L��5��y��-t!����``��<C�d��ͦ��(��}�J�~������ܩ��S���j���#�"������f��/�'+P�^����(Z�`�5��_ԕ��y3�(��8���.xA���f���f�ƨ%!)|S���?��x��~�|�H��r8�'#k'Q��}\����e��O~���ku6P8zq�h0���.��e��`�ȭ�;��R:Tڟ��#3;���Λ��œ���Q��E$���1ಘ�&SKq'�֍@iM�>s��_�cbiI�A0��%	��F=��JI���;@���0 �<���s�<ʫd�iq�h����z��� ���O<�M>}H�Z��ͅ4��R��7X�m�OC*�B����b�c�,=3�]���Lޙɓ6�s������2jh�QZ�*�G2U�zY�J<ژ���b��I��߉��6;��d���|�C�I0�|�ohI�Ȏ\x8��0�oLSB�t�w?/'���������A��@aNU��<�|"��m�`����]؆Q!�g�h�

��6�̩�OS�w������*�F�C��Ƒ:5�(k�u�{�C#Q�g�tA�|��"LMo^����a�7�8A�B���X�v�Eޒ��p9�e���xļ�]�)�yaO�����*&l��Sk�c�K����)�KMU�2<*�����Fv�7�/y?j3#yT���F�IX)XMIs��C�9w�\z�/�_��O��7A��
���Q+ �	�v_���0D�BQ(F�c>_��R���$����֒L�A����-������H2̠��(r�!�0�����*�2@+�ȟ�&�xR��	D���n���X̦�c���H��yh��?>��]��hKfLp�,�I�g(;�q��4��#��a��x~8���N14Y��������0�h@����<w��*۫���UXG;��w�ak�}[�p����)5�v��R�zFFFrK�
�p��HJ�I���<Iڣ�̈́���GGG�cd�DG<�	�\"�Y �@���#E����b�~�:�<�6!+���Xi��477��6��/Ό�L�lT�����(�|C@N��2���M�P�{�$  �Z�ra���2$(ŏ}ļʦf&����G��#�����7���G�v��0��1�]i�	�Ϝ������q��Lv!�o۱b���I�xTxCm�����bxZ�=�	 �h��3������v�d�+�Y���²�����9zh�(Sa�J��RPZϬ�45�˂Kκ�Y�A_ xDlST��B�r�Q0jjj��������5��FX4ĸBWq}�W�gm��[$w����U06�eƨ[�;��7�yR8J��fP؆z�dcK�vc	Oލ�������_^�����f�E,�DE�2��8�ũ8w�ʝ��Cʅ��F+T��|������뗮p�9<pw��y����4MA���vl a�*b��1�gȚ5���!�M@@���	��-ë�������?~b"��ЮҰR�;��o�o���^;0��F����'�m�
Z�ہ�@T�Ә3�+U�v:e;�FO�B�Y�ѽY��/9n�m�.(�yo���:�j,9�Ơ{:�w�.EN�t��?�J�&Z.�� ��\	{%����r�|�p9���&+��d��3�B0{��Ҟ�H��q�f��P���`�����Br}MH�R�οh�3����%C#g���HM����
���g4z��=0���%]ŋ�$��	��&`�˕ٵ3���)�*he
��L[��1��*��i��B�� �#hq��з� �í�^9��)�XO�U�<��9��O5@<�J�6�k�VW\���8ʅ��*��b��dWX�6CJ~���[ב�6/����3dv��ɟ����n{3�4my۞��}����2���ɼ�^!2<�3�V�kpu<+l%)L)M�Q��)u�wX�Y�g�t5���,����	]��|$L6~�Ys��rA+��R2h�E"NU�Poܐ#�~�h�����I�e8���9�L���\��`$�@6���#�b��W��Z����JĀ������DŀQȘ�*Z���ɢ�,s��U��ب%�3�L#�Ή u9���a$^8*jB�@Z`m�Rȓ.���A,�SN���_p�8���@���Mʰ�D.w�/W0)�8��ER�8���>:�6�Q�D�(΍���$�`�\�\]c��?+��L
�/�e{��ƕ���Mo���V6Z��&6a�L�z��X�Y&��_��c��<�؄�O�;pD�ԥ~VӢy�S";B�6���Aƹf�Zǃ�h�<3�ʓ�G�eU;�e�:����c�˲3f��_�5�����#�]GTNҠ����ӊ{�[+�-�����a)����zF�qь�l�Ro�(XBy �띓!��-%��}`�;?1}�43f�9�0;}�Xl�d��!cd5�?�-
M�pCi��F�7?�u�Eo�S�H��p̡/o�Az��*\�$�E��a��m����L�֒�P�2���D�i�š��x��w(=�N�~5��b�ehp A�e��'�v��T��#�~c�W(�BC�3�G����`�2���Vzj3T'6������ۖ��gal��q7Ui8.\��J���$tH`�H�j���
S����T������I����BZ��ُd|]�eŅA�L J�0k���Xf���6CG�S�A� �{�+**�]M�AR|Z!k�Y f�!��Kx�#�#��e�Jd�{6��yKa�> `BC^.%ԛv"�YNg�L�1�my��CIE+a�]Y��䘅ܴ
�z�3�p���-8up�]�E�?������/.���$�F�/�:1ãJl�R�}�U�"�s^,f����_�}pޔy�A~$������ps�Q�
9�!�9G)���b�b���*�g�e5;e*�G�����h���fq�2C�U��Z�H��Ľ]����|�7������~�x�u&���,��  z� R6u�âK����EA#ԫN%^2Nj �Bba<? �C�(�"�����;EC^r},:e�떦��Yv��o���\={�C�-Q/}�-� �m�"����+ACCN�jɡ��Q����`C�-nm1��)Ԋ'cZ#���Rp�c�}ZR�����F���Vj�ML�����!�RW}S���rd�<��C,�%UU�oWm;i�Oj��g�T�I��,�&�%���O����	WR��bȫ@����v�� h��F`�N�s�Z�o�Ѧ˜�t]�0� 1�|:dm`�dE�.)|�J4�o�U��@%�Mg��)K�Aʥ%�^�TJ���م����ƈ��È�P#���r�q��N�/a�*7ʦ@H��:�dƂ�Ӿ8p:�m���<�Nc~���\~,ԑG\������W�B��׹��bV^dƌo[�qHw�l5���m�qg)d�ʓ�چ�v&�u|}V��Xu���w��t6W�~��~�9D���q�H��"0y��]"s�[@�Դ���5Z�K<=+N�:)Sh��`�cf�b�3�(
.�E�TxD�\�'�n�0�o�2l�s���*PfS�ހ}����-�d�K� �}Sd�D4zUG�JN5U�l�]"}�+++ˏ���j�_��d��s�~�c�'R����y�0��u?�B<�_�ur̞j���7;��4��%�`*��n��3l��d��'䒌�q!L'ڙ	-��{?S�ј��_߯�q�he��@��m,U3�:�.̸��q�o(������\�������	RQ���������~�Y��<OH��c��8M�`��Vm��`c�Z�����{��׃xsqޑ�W�}L&��*=��:H�!~��	Ij� ,��H4=K�W�|[�֙�p,6��Sea�`�ܣ$�x8K2��19;��Ty�,۳bP��W���_k����E>��8 Kl�/��,�}9�xhw��K�S����5�W, N�`rT,�"v�ь�O�M�����=��n�z��"�T�MY��AuMw(����,v,�^��.V��q:�~���������M�YY��"͢��G/sm:Md�M%�d4�̿ly�#�ӛ\'�8����0�r.V�W�Qa3(S�U�Ck"�t�����iY~� ���c�:=�>���n�
8��@K�'����ck�k�~j'�d��r��+�OA�>v�K�����qR�k�1��(H����yZ��A�KR�z�o�P�t0��z��U��s��$mv<�AXg)�s��U���� ^�ؾ:h�/�REJs�����
��t�n�����zV��7��U���9i��_�����vm$�	��S�	�˧"�{.; ��`	�̈x����dn��0a4c����w[gb�����b�~�qq�����4F"v��H.f_�0���1 E���V�aמ	�,�����tZ\^Ǆ�2�RbYS��@}�s����~Mz{8�#�ͥC��k������&�9' QRUm
�����}�(L4No���CV�m��J��#���RL <����������Y[��#|Xlmm-M�R�5�i�����n�nov
G��$	�6��ܝɀ��̏�w���Y��#3WHu���l��qUN��Y�?��DH��HF��ҘI2��b�D�6�;��T���j�w۹��6�S	�E��f��,�.H!�AI3�58a�^��#3��#�:�w�	��d�s{� O!�����$Jr;t]q:!^�6Jx
;��b�L�L�%��@��Q#I�)&���H�����j��Nޙ?��6�����8>u]��GyG%=�s�\#�P�uݡn���?�'7�,�ҙ�������%�Xg�@��7��ߑ�0kᧄҁI��?��|~����(GD��\��뷽'�;�C1h��	�?��mSm�{�/�|2��?���^S��p1pþz�6p��/�?L4[[d���g�5�>��_�F�BO�^��poH��!�Xr#p�y���R��D�2���݇�)4���2�f��gӷφėH��	&:��D�ѻ�a�~�dn�ì�|�i�tK��|4��q���	ߵ�K��Иd3D�dvLTVI�XxU��y�|�E�n��W��%����P�J.���&���e$'�Ax L��q��9�!8Sݟ�ʣ �ui�%���xbP`Pg���=u|��cB����ez$��M����u�rs�yDȡ�0��.��'XSn�?c7^&s�D
�y��nAC�Ώ������ɋd$m��_ڪ�w� �W$�" c���M�Zyu��>�+�U���҇���br-�u���dn�F/�͜�6JHo�Tn|�~c��{DZt�[k$Y�v�"�
$�o��z���`��P
�
��!L�]��ǥ��
\
Z�,KU��O�0*�ț -��
�L0#w��{tx�:Dlʓ�����|Ej���:�'Ü9�w��\Ms�ÝP�R�B�M�#C����խ(C2\���hyȟ%_��<~�R]�Q��|�g�0�n���u���<X"=v�v1�;�@��ú�~`>4,�u��>.'H�6E ��#̭읞ka�)��XpQב�)����>?�[�c����?dV�9f,���۷ǸMCX�{�a�}x���В��� l��Pj��Q�٥�,"d;��Ls�'�V�~ڰ�S�gV��LK������Sq����u��vGL���L:�.B;���Gr���9�z0I�CR�J��3`���5��ߌ��D�*,�0=���g^e#{�$uCe[�_E�^I$��4á��Y��8�&��4$����.R�bI�����+rӣ�w3���m�ߪ���}�/�IDG#����m�;�bQ��9��|x�#��F�}��!1&f����%���#j��Gw��V��WEf2%Ś�[$����	-�x�+��U8��|����>eC\�o���-�:❐�6KRxQG܁H���++Q�]��V'���������	6���((R��S��ֆC�6v����6(�0�"��������I֕g��fmk���N�$/�O�e���n*�M� �"8NNZ��D�~�>*hPxq�.�|�DY�m�F6�������N��X��I�8�!��nC �81�U�W@ET�f����ς�^�J}�(ci�L�[u)�X�k^�z�C��+�9p$�<�[9TU��<�Ue�8�1^���X�vV�������Z�t���4�����X�.}%A�aC����5�<�ܽ�"@��#D�'����ޫ̎�WM�n�b��Y�k�A�bZC�F>���1xZiA�/���'$�;��-����=�t��n5���[�HU")��U�'-��^5�"y�r�v���0JŨ�u�/כ$��'��[zP���p���6��_����&ωؾ��g�g�܇�����i�Մ��X�']�Z�α+������OᢺL%��0��0�sE��]UhlM�8ac�%�@�!��0u�Wj����׎O�ڪ̥t��������ͅ�\���<�q]-���i1��燉��4���	�)�6�"��6�V`~ڧ��s���y��SA�*�tq�S	�8у�0�Ⓥ�q�q�=S�[�ё+�T̂��!1t��(0��F�	�����B	#�Y�<����N�ҵ���3�'�Ί:뻲�9�=��1!�^Ab=c��Ī�JR��p��+5�x�P1\�؉x�p���
��q��`���BHh��'e%�A�Uj�mK�|�	sէ������g��z+��%L���گ�� �έ-�VMڷs��G�M4S�/�g�Be�tZ�3�����&����}hQ��t�2�.@*;~�W����F�j�|	3��UaGU&����dm*��F�VsfI�3:�Ր�Unw\��WG�vb�n�7ZiY1�q/�_�����[�Ћ���C��0t
J$+4����{�d`�J�歘3�$�`B5���9�j`�/tR9��wNk��^ �tVzCWj�ܺ��V�2����u����d��?��y˼�Qf^s�ꙋ��ʖ&����I0�����yK��"⬓��G��G�B)���F�J[?M�&
��D��|�4G]Da�����3sG3�/�H&���Sh`�#B�Q׶�ɡ=�I8����;���!B�fde(j��LO��������	4�2��i�S��2&֖[�{P�����=y�*!tc�a<�Q�����B���p~���*ε�ܑ]�O���A�=躻�*JB�Vp�y0��a�H�ag�o*d�uB8�FfU�5�匐��9)�_?<�Rs�&�O�UR���r�ט-4��@w�I8�9ܳ�IZ���B���<t��ͻwU�{"���$�+�o0B�c�Ā'.`#�a��h�f۷�>S���3�d֨�{S���A�v�=��[;N�u�D6�7'�.��~��)q&��	0T��U� h'�*V������m��ٲ����2���4��!B]*���Z6�gD�>�bGL8v��ް�tP��G���)��[���N�+p�U#��j$G��{J=��.�[5�i!0ѓ)ˉ}AQoK����o�l�ۣ&�c�o#���w�����f��� �n3�]^�n1
S4R̕bz�P�w/f
�P{��i�vfZl���F�)R^dnb���̩�zO�Zk2�
W� =�4<�	y�d�}�O��Tm�W������𦶼���A��m5JH[��/5��'����H�+L�3���9=a���U�-�^G��C��γ�5��$�6�pl��Eda��A�N�F��j��ӝ<�𭺑E$DAlwyoL�]Ӹ�"8'q0Id�+��\�����Q�CQEt�\i/m�p+�e�,�Q��*k���_Ȓ <����|}Iu����R{or��!����J��g�c�h�>S�e|�O��Q(<��R̽D��zL��H�nۅڱ�2�t�LX;�%?Q���'�R�m{ˆ\<I|q����wl���v�о4y�'f��v9� i_ս��ƀ��Nٜ2����p,�SkL��x~�5T*/�hq��ټ �T*kT67����#��������V���[��l��bN�)���#FQ�8�O@�ֲ0�`�+��Y,��X� //V��/$����{6�~h��j�}4�l�A�t�7�T��`Ug��ZXҤ��H)�h%�5m�tI��v��ƞ�0[@��n��ބ�$�^��,,�ǲ`S��~�t�z��!y?�X��⽩���GU.�R��&��h������4���=��=���.���.S�[dr���@˗��m�\ʱ�[t`�e=fPl_�����d���G���S���#�~P�D���ݻ��%?�L6�����9���q���׵�e��(��j�`�|�:XUNLf����.�/����|CĮ��ვ/��;�L����N ��%�V��f5G�Q�x�;~sV��
�i�[$��r1?���ߗ�����0�K@ް`D�ϔ������ ��WR�zb��;���*�c��Ъ(p���t��܈D�Y�����)G��<�,�=�B�j�ӘыBk����(�>UR�O&�8v�%z�F�N]up�)��]�΢ń*7�J���\���J��ԴI����'n�s�)�_�D�
s�3��C�#��;UU�rI*��庘���q��4� ���^����U|��W�-�co�@��)c��-�G�¡bgE�<��D�ʫ:!\7`$�$�S���ȋ`101asA���}�(�A��n
�5�6��J�S�Od��ak�su��d�]	1�]�%~�b�+F�zJZkߧQ���z��&�lM�>+>v'�������݀K������S�[��5>5s���o1�ʦ��}w��aѳ��o*)��G�!�]e�"�<�]U�� %[NJ��/�\*�?����|��ן���IC�&�&���+;�����C��w��@-����-�.���:")�R��������9��Gtw #����9jH�c'�� ��Ic5�Ve���/]z�xP�9s��P,�%����F��/>H��P�3_�܁�����s���B��l��ˇE��{�ŃgdW��F�S��=g������S���y�X�z�И.���d�N([���SYt�#�˺�ӥ��æ�w%H�j��-(�[�-b���oZG�oE�iYf�3��18�� �MYN_.�P��%��{g���=����қ�21���O>�J��)�׆��;�z̲�Mp)��f}u�ݸn����ic��A����y�e��}� Z  ��F�����A��S�t�l�}���ч���iD cm~�5_?{�/���R-3,hQP�ĥ�`S]�E�GjGk����R�7ӎ&˷��O�P��}& |3 ����]T�5t�^<V�x�J�sh��}�ߕ�@�I_\��	J>'��I8�ͬ���i�T�:t��9��GO��ad���������Uָ�x�%�P�gd�We��-���&�����E�H)f[U��<�8�T�`�Y�V�Y����C*��eΈ^S�� �SuLȓ�������c��2=�O�G�����Ds������؉c�5�����Qq����גa}�-�"��1��V`UXQ{,�M�WO�����:'e��#�.Z,8��C�~�5��<-�E}�S�Jdy�J#��<��d-��M���23#""�F�(U�dU�5�t�y�$(l�5k��>�[�1W2GQ��	���[D���}�7�R�0b]�՜"�D�;�rH�a���A�$�ᮓ���&MV@� [����{�I�eƺ��A�i��W8���<:�������חB
���r�	�*2˖��L���.X��	��8������Ñ�F�I�ҥ��q��G��a��A�Ѫ�,Gu�}��	�,-F��'
�ň`�6�/WTD=[o'[�x��U� &����vN���A�D��AՇ��f�J�f$�y��?���yj�I���Q�C�p���̒Z��4d�B�I�	�r�zo���i��u��̺�R������R1���>�9��N��Q̰�h/`��\��-c��E�,_�� �YRp	��8���84T�_�Z����`�w��&\���B	��ޯ����<a5�/^����Nka�i���[�aI��b�@}%\đH�7 �݇7L(	Ne-����e�o� �XvUu/�~�_��'}
xc',����y��Xb�4�b���U�Q�}���B�4�Ѐ��.�?s6Wu�scg�97e�O2�;�g!�!9�5�ɿD�&��H���Ҡ�N�����R�m��8b��*Ӣ#�,����[	�cA���J��O��oއd��f��]M˥ sۑ.�-��Pq7��e
Y����H���w���3������?ۅ`�`f�5��o��Ҙ ��#�J�}�ďS�$�I�(�F�e'Y.m�̲�r�t2#v7J�eivC!Cz�0RHd���Ch�
%C�Ǉ ���K�O*ҕ�79!��A�聢9w���))i�0 ��^�$�gxQ{��h����zoC�
fx�9*r���t	&�`��܏]�W_��a�m���4��*k=���Q1�aC+	�Pw�{�ӎq�֍��Q*z{���D3�������W�-��Jatjs	�k����Fs�Md���߁a$>"D��&�@L'��;����"���	�����	�%��C)vsC|X����S�O	25��>A������D���"%ty@:��*�k���|��J��?�yw�;ײ��O�jǵl�@����w���Y�c�y���,fV�����}
:w���<B6ꤠ�����3�T�l�ЊB�N:*P��;5����C���������D'B^�.�ȕ����8L�Y��V���S�����$2����N�溳��q&u痭�}��MƢ�ifS>J�����ٞQ�w�w���t�^{cߥs��tk����$���
���@�ǈ����x�b�Y����1厖�>q�Q�I�AG��RQv�o�p�J���$��F'v��W#5�\#s����	e�"�f*�r	�K�tsӐ�>�����V��H�HT����^T��_Rps���f��J-��IB�qtAkiWtnD�_��UG�N��4��F�z��H---��	��秧Jy�44#�E%�q�ဘ���)8}:�|� ��(������\�ϙ��[�q�SdJB�P��V�-�p���G_<;,����F�$�X�i����_̊�����j��L�eu1��"Z�J��zX��¼z��#�xhMl��8Z٣d�Rhe����d҃�!�� (���ؖ�����Z1|�kh�,��-ZzF{̸���h�$h�-��/ۮ����N�G�-���r�
�
hJ5����� �I�e+�6��7)��2�Dy�B֞���!��'x�:�+-�$��fG���O	(����y��A;^���ޘ)��K;|�����33�����V-2��<����_O�-J5P2��4.�ł<n[l<8b�bK�Y����$/�E7?�|��%�*��Iђ�P3w��1�l�X\���IqK��w$.u����B��3[b�!���{�-��)Nv�fs�9��|&�%�8�C&ŋ�?���W{���3�\��:gx;��%۩��g�����{��p5���I����t �Ƌ���������vQ2�I�_��Ì�/�����Cj�o���*�j����6��Q�Z��(4��)�4�����6���:��>�]��؏s2j<��FEH��&�b�i-f#�B�С����PU]�^�x!|�ܵE6F�y{1yq:�BXBg����1S�#߆�ף�����K4��%>�DS�h�uЙ��ig r�W
G �<����
���_��!\�j�ۗ%�hrɧx� kk�� �jjw{�"�7%ߦ��C3�Eh��t�=���c�O��s�-p��u�m����Y����,����Ø"��6F&S�Wk���JbR]��|��Dm�!�N���ַ��BJ�����L@;�Y�fJ���ӆ����|]��-���k\�f(�]&�*Zy�8�]���*�uȫ����"Ő�K`}쵯�AAYJ�8�NLSz�'��B��U������ގ�U�-$o�rFWY�O5-?�F�c���n���?��ֶ2��%|���w�`�z�<�^�)V�.2�L�/�ѻ�w=�����pZ@{�<�<�깉���R��x�2���i�Z;�I;Y�m9_2��F;���3��,��=;��_Nϐ�5���>��]As9�ٽ\N��+{6!C�_��3٫m4$��;�>3�zw���C�Em.mծ��QB��Y�-v��`*<l�����n|�>����Z�n�����d`y���|�{�t��O��0��W�f����gc���\H��Ha���F,n4~��]/_?AQ�o!�'ʠT������7}t���~n���mkd��	���cʠ�Y����C1stS�rG\�k�^�J���.�5?�@DE�dp(��muF%����N�
�$�GWr��B�Be;V��D��Z�G'�7���ʑ�;ל���b�녻ùW:$��EJ�P&J5���ZYBK�Of����|�����$K���!I�t>�|L�Am���3���5i�)� e�sy�|a�a_�W����ۗ��V�ԝ#�c���� �O�:�r<�n���A�n-���8ؽ���{��K.NOy���V�kǸ��r�95��V5@W���Z�\�w�gE��
2�A�#�>���o'�#&ʸ@��k�T���TUe4��ʚ��3����(��@'3�FT��MG�"��"�^�!o��I���0
.�`�	j��"����Vk���,1�4T\G���

>�7L��[*�
�U��ڱY���Q�>�$?g`^N�f���a-(�5��3[3���s��u>�ܖ�^�u>g�[�|�ha;mϻ:^^@����j���$�Z�z�BB��sħB{�H�D��/�?��ä�{4�K�k�^*��j�c�U�;��JN
/��@�|I!�G��k�����^Pg��s�L�?nO�抂M�8^�����9��eW{[4�bS�nf��e���C�ҵ������~I��7e�����\a���x,���,o>c�뿑\'��N�a,�#Ek�|mN�R�'j)��M�Un�� ���:���m���ۍ%��q=�%�����g��L����� ۙ��o������`R�5TL����O��f+��`��������tA�T�Y��y�����X=��mm�]l���>�/{�_1��i����	��Pk�z	y���kϓ����瞓V44�y|�a�5ק�)�ĢLމ~��僬��ӓ���ˡ�� r`��
Д��b6��y�q5�������"721���F�&������n��C��޺Ӕ��Hk�-%r���/���/o�9B����16K�[v�~�}�
SȥY!�g��Yd�Z�r3�5ⶪ.O)��m��dt��>���@"�Ef�);s��쌛�m]:��qRZJ�8L����I7*%yc���m�0W6�u��9�&�⺙�����31�^��%`˘!�J�Pϵ����4mx���+%}�����υ_iR����,�|����C��L+�c��_fʃ�|���5�w1Q�X�ö��P7^�}�<���G���@�T����c�묻/��>��O�������7��g=�� �>��7��6��931�v}��>#��ar�c!k��nW�c*��yG�<^�637Í��}�'>U5Vb�Xc O�Ҿ��`:�$����[u�s�Y���(��u����߱PP}�%�B�,X���~"�n�cZ�yb��7Uޕ��q~.ϿŧzmG��Ƃ\�]��z��T5Ā��mBo���d�ua��t�h��ʹ�(܀|�?wa��&,6a���H�m�u�ߴ_�S�֊S��{X\=�\3]�
8�<=������^�,7pɋ���� V(M�E� :�:Cz�x��+=J@��@� �maF��̥������5g4p�D1'��f[r����x����P���v���5a�~��<]&�絠O��_=���z�+���������Q�!A[ڥأ��;6���D@{*d��Ĥ`�6-\��������_�t�kn�����
���.[e��Y�Pf!]e;q�Y����;dtV��Y�9{�r�	Q2��e�p����}�������������EXT������2T����aZ9Jf 1���S��R��+��n�Nk�es��:�A��A�־��ĂP��tL������|��N�(�̸r��,�`nf��m��q�%����} �M6ϫ�n��[�{��eH���u\]�����]�@�S��^-��ʣٍ-N�wv}�R��Ƈ�Fꈟ�t2��+G�~5�����)��lWcsm�i-������,>'��t~����2���ta�i^�a-��XO�)�c�]{=�c&$�*ݢ�O#lĞ_82���E�KV�e
��u��}	T�y݅�2�u}�q���{�9�r�Pa���{��x/�c�wH��ַe<��̭*���%�-�w���/?�,W �O�9����߳��K?\� Y�[KM[5�Ty���C��¨�Vs���l�~��E�<�}���~{����~S	>6���G�VUŶB��N�&�lh2;��دHi�����!�-)�f�����n���Q0w�(�z����FZ;�����QD��Я�z[��H9����a��'��e���K��	L�G��{�g��)B	�;�0_iF4�(�ab�'�B�9W]~Js�����x��]B����t���1tH%Z��}��eq/�;��Uc
jW���Dd���R��<N�c.�,���s��P8��-v;/��1�
l뿨� �Ok���ܬ?���ޕ�>�	q���G_�4͎|�ѷ��7�*5x>��?V'��/�8��5��<st�.��*]��Rr�~��������<�Z������L^h�.i�<��F�@ m8mr0�kn���̝���B93��Ks���_�~T-s��sj)I�M��s�3�y��9�Q��V�\��=G������D�Gt2�Պd.ǭ\GT��M�6K�fT멭x�mTx-��/@�2�ظ��0R^�T�zr�Ѵ+/6��*TЇ���R��"�X�݋�ẖ&���G��Jj�)��X���;b� ^�ؾ1c�=F�#��W�D��tH���w0��4����l�Q�#�^���̾.�_��p�z0�O<ϧ"�����B�׋�3猭�N�V�{�ac�uF�z׳���X9�Uf���.S{^��aDR�;.��O��i%ϴɋ(�	o���{�~�-���룳%A��%��&�=���վ��N{���~�:d����yd�)�*��mĥe��k��rz�~S?߉���V�?�P[z푖�ˁ �i�2�o���PY~L�1O�;�8Ja�����4Lw����/�t���[cɐ��5>�'�b�z��!�#k��Ƒ�`��#��
���¶	�[D���}�� �S�O;�f�E�k�I�2i��1kJ��W��0'%r�	�%���Z4p5jH���?ЇLe4����ic����.\s����ՂZ)I'�j�1�Ws!�fbKTJΥ{
�7r��{���X�o�v9�~�]p��.
-c�׎3M���Uٳ��eg�ϸD+���'�ٚ�,)���ɧG��+3zxHD�j��IOj�\�tR�<����L]Kc#�
��I����o�.�E���b�c.jm!V�� �K�[x�F%g� t��V�Ja�����?&���ȯY�Ώc���O�M!��B���(
.���L
ț������n-+Η��C�f�O)5֘��Ԋ$�����B���X�qe&!��X)t�����m=Kh�7�'~S"�,��Q�9����^5q���Z���!w����S�4,̅,^h�uE�8�~<%1E��҂��R����R\2���ZEL9������7�K��r�w�6F���5���8�C�6c5 F���9� F�,����ZW�}`���VUU�;�	�):�ހJ����9��i���M?p P�y$�
�O�^y�����y��#��"�x@E��`�D�U��ȯ,�L��]i���h8�p���g�DWYR\�-l��p����|��oh���&�Xs�QL-�4z�W�[hM�J�0◢�{��g:O������e]d%&�\W{6.�_�!L��;��g�� Yc�J叉�4�;�4؋d-2��i�͐�ng�9��XO�H�W���mZ�Ŝ��$�0/2z1Ñ7�T<�k��M��t��k��dR��ٱ���U�е�L^s����Lf���F����U
G����rɜ��^�A�2��{4�ps]����~����l�ᷱ����߹�������[zA�u<�)B���֮���'z圛�97�Z$���/:W���������0e�&�DN|�����_l(vt�+(�U!���^������{��Zz���¯��o�c�F��q���;i*�O�"� �z{�Q~�}?Y�������	��]U�|ņ�jpȫ�����º���&��Fތ{�@�,C��۱��͔�G������Z�c�	$����D�C}}��U�ph�ִ�P��q-T|T�^ԧ|���B�w9e�;�\��U�H:;�1�닧2-���է���q�K�2�nnO�����PoS�3�P��Y�D�vp��-n������v���Z��DSQ�8e �`�G�^
�}�nt�>o�+��Y� )Sz��;ar�#	�ݸUnHs�4�uڧ��ᏟIs��N�/	C��r&:"]���)��Lй!*wQ���*���\|B�O�<vd|���r�d9ܤ�1��"Wz���eXh�����˓YY*��Y%c�M�=��:?�ȏks�{LI�%f���W��G/D|�q��+B��C&�ך� Nj�_Sb�+�
.HS+&�T.��Tb�(��
�5ns�ν��%�>u��ܸQ�8�8�r½���^߭6N�k|N�މ�m��B��Fz\Q��צ(a�%�GPV{A1��2O���s���
p�i{�)�9	{��8.R�x����.���;�m�nV� ߑ�
`��1m��]����YZ!�@L��ݬX"�5b��V!�H��!����"��`]s�#	7�<8ٴ���?<Agۓ�w��lkA���Ag���i�Ǫ��D���+d/խ�����*L��%@�v�p��qA�_�t���5m��PK   ��dX����H   C   /   images/8e6e9996-4250-48fd-a42c-980e5b13088a.pngC �߉PNG

   IHDR   d   4   |l��   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��|yx����=[2�=dOHB6H���Ȧ�
����R��jk{�t���zi۷������R�*b�V@TY!@����=��d��=�L&$di����I~�[���g��9Ϡ�Y�����b�x�Ǉ���'NwC�R�j.�s��u�B��Z�?q�'-jJj��c��c¡�v9�v�w,��G�O{5:L�	}xߋ�mgI34�o��RB��h-��%C����v��:as�q5��Q89O�2{{Z|؟����,{r��
�:6B�U������B̞1}�������N���*�Z��Mya�������\.}2��Á��V��P+ZL�o5M`�����3�)++3(o۾� ={�ɖ�j,tOrL�_�:��E�]�����������S�qy��Mʰ:7�-Σ	��my.�cA�	Ĭ��Q�Oar�e^�3<C��Y�e��w���k�5|���Pw-��X�'V翐�����mGOgZ�.��e����@�� B�@t�Q�֪eR6��f�賸au)}~\���e��^\���RM�����FNz2�:��i'���G���E+�AH �F�9D��59�X��5;e��DJ�V*����8~z�ɷ&'�{%8P�����V6w@�V*���j4t<5!6�ʖ^�4t�	Wx\HU� c�MN����H��BhH04�h��h�Z��׏��v�jơ�N�t�`�0|=0,�H�����c0(*�I�t@���p{!���1==�s�0-k<�b���@Q@���fC���ӭ�8^݂/��Q�a�٥5�"96�/k���7O�}s[��*��,�AV豿��������7�"�X[�������i!��T�wAI㓑7m*V,�A�ށ�GK�i%���p��Ac������D�.h�k�W�I����~�(��f�c�iț<������zss�`�utuu�HI����k���U���� �m���Q�D������*�
n��Wb�j�3�
��	hii��`�
!�������T���a���������CxsW��c��'�e�A�ų"`�*Fŧ�jZpOON�����W"V>/y�%!xx��#8�h)���D{{;��܌��^!:�����0aRRRI�187%%a��|��{��8��.�O��9��zΚ��-�I6���+������������ݻ�u�V�<yR�Ɏ�d�J�PZHFF�.]�U�V!++	I����k�?�8�����e�U�5Rg�w7Y�ƣ��	�"'#���?�>���
M&�yY�F�҅�����~I��r~pЌ#G�࣏>�W_}%��K��S	�������E��zsss1.:wݴy�����wa{�����I�ya0R¼x��B,_�� X�"�oߎW_}� 5�e��F=:G��Y,�8q���X�~=��<��Cb=�����"�����r�Pغ�f^��һ1))ڀK�C����}&|Yg@u�Opc#X��S7��{�,CHX�X;�?�	��n���3�*��+��y}�x���
Q�w�yG@�я~���Lg*��X$��ފGڅ���9���T<YƳ�Q��Y"q�������q�F�8�d�PrK� MVE���dF?i�iP����_��_�w���ϟ�I�&�?P��ڇ�]k�83g-2���Rf���$���g)�C.L�g�ñ�%y�B4�9ߣvS�䖟X���X)q�l6�7���/��Ʉ Zg�&�ؙ��
^/���t�J�`��[��o�>��7��ʕ+����_~�k�-��q6&�&�f���ibFSS~������iub��� L�LG�����F&Ǉ�h���@{[�O���|�V�Eyy9x����X�b2H{��ף�孨��H�c0��`4ۄy�"#)
��:8u�A+ٍ͋9�0c�x�t�CK|>6"�m��n��¼t4wP\݊�-2�G�����߂x�n�Y8��r��100�g�y���D��`�൦f�#�,��(��C`��Bz��q���vY�^�Ǐ�cqs=� b���Խˡ7��%6ӛ
�(f\+��������i30uz��G1�?%��9-@�]\,�f��T)�ع��� �F#�q����Ǵi����v<��ð�Ւf���z�"��ff�AO���!� ���us�VbޔT��eAv2��}�
'cJZJj�x`�l�,vܺx�\s��E��?�Q���o]���q��>��h7��C��&�!o�L�Q�~v��1�x ���D\�R���܂S�J`"p���{N�����GJ�<~�BԾ����HLF��G*��U� <"2;v/~0xL��M$���?�ȄU�O9����Y�/Qdm�������(!�_�BX���������n�K�Y�y�t2o/lD���l�l[��SR����퇫�EI
rRĪq�dQZa0�SSq����Z�;<XK�ha�9d^��5��ƙ4�	���� Afdgaz�,YӅT�����dM�QQ(:p]�bM,K&9�/F��<ܽ��o�aG|�y�z�Ǎ��fbJN���mۆM�6[��=u
M�-�����u ��i���iBPp%N��I#<����7^}�>�P��^HB(������=�P0W�jw���G���0g��N
�UL{�	�����ാs&���6��d塺@Y���:|t����Š�!�E����)QX4o�ģS�Nᥗ^b�H����s|5�`��
�u�'H�3���%2��x!����=��)S� �<����`��F�u��s�a@8�'�����>�'6,(�C�I���IS'K��+X�J�H۬V�\32�
$���<AC~ۋd���q;�|��K��c�	|7�p�fcav�QL�B};�,Y�6�-���pk5h�6�bs�����(�m��RJ�0�,�&�<��M[(����u�`�,C���f�x1��^{}}}$�-��ř��ȝn�:���!�ޡШ��{Y�V���B��OwJLe��Ĉ�����3SQ�I�0À���ɈFf��{׮]�Y[8�O�1]bSvO+�&8�%��vv��7�L>�4-��$��T,�����g���Ѽ6��P޲���֓� ���LEc��fsbDPf+9R�$����Ҙ���51|o߀e�^!I:̜�-��4~�Ν�r)S��|!*~ː�@8]kHl!�TС$r��x�?b\$&Q��x�����vYI�����{��c�Q}���B�<2����l��ux|�NԖՊ���\��`�X�� �W�J@#Ka��Қ3o.N/����~]]�$Ry�iH
/BC����$^�)J���tW94'���G�+Z׬�����?���az�������n��p�.X��;�e����jQ���Z	�LKANB�֛I�J l�Q:%rғ��B�؟2�<A~�
[�m�B�g���_�j����3y���db$��u��=zT ���AV\��p�5��C�ʃ܌DZ_ �/��R\1��#צ䎥�u1��3� �:>�aוH�My�S�$�˗/��w���}>�bB4�����\��:O��:�؂�'Iʔ��-�27���ޞ^�EF�ű��H21���Zy?+ ��MYc�WjpHP"5!F��K�O�<)w`e.���\�^��5)\^���K�Gme����Sl���'FQ���k��R�@}ȣ��U\	�I����Sc�p�e�����5(�
����v��V�K<A.Nr�NK~;n\���Tx�еJD���ߜk��b�j��Q��� W
�m���?}����}��a �{�A�/TK=����%�`���ݗ��QA���6��5�`.E(����X	t�@J��[׉����!-�r�w�}�af5�!����u��Ā��:8V���rrhw�`YBۆ�����-�@��O�Juق��:���pY��D����|_�0z� p9}�Kz��{����0 V
B,,h�����5ea-%��;i�<h|��XK�W�9�:����؛�{����8씧8�\���������/!��'��i�)��}���X9q1��N�P_�jw�)��Ff�qXOLL���o0צ���M�R��C��;)	�Sk~'�D�tW��p|%��D����c6L}�UV�v��a�U�*�4�r��^�N�db�M.ޚ-�=Oo�	z>��D��ϻMNt�(�NEzz:"�]q,��%ם8��=�)����b�F��Q¦PKi�=�շ����p�qM�,\��O6�=h�����ڒ(q�0V�F~���+>�
	̸��� ��2q����;?��w�."8��}p�)��B��Yݨi�cf�4����P6�EEF���q��#�&�G�'�����)��mX`���K��]�b���={�\�Mϭ�0�J��݃�is)P~�+Ic�����L���66 ��U��O%�����
�`W�J����A��FC*�{x����%��l�����cٲeؿ��.q.\ ~����,#-3�Cp�|��٘��.�x�:�a�:�;l�-s� ;;��@Em#�\���"�c�� &6Nji����F�]u8y	�q|��[Ɍ�uaP���rD��$���5��g���Ȁ�hjmC��$uAëf����Pd�p����E*��z=v~�V�^��d)D�R3ӥc&�+Ŷ��S���N>��gS���r
g����K��j1c��Z��\Y<�&V�6���:,��EAA�Ν+JȊT^r
�/
���J�Z��ű�<W9X�آ��J��bs��Sb�L�V�^����1v��
mnz�Y�E��6�����Id��3�>� ~��_I�ݻ{�⑛7��Cu����}Z#�`4�IBg�Х�D����<!+e��Ipsб`��N���{�;G5�.u\l�$nڦ�����;3O�G��?���Ue����c�C�x).(�P�������ix,�_�B+[���>�2��6l/��-QC���C��6��wO#3+w�y����U�-��$�͞�#����W��9Fh�>6�4�Y��Ox���C�슷�<���B���Al�u�F�9E�1�s=�� V�E�z��'۱�D��?Gv��{��K�PY�I!.ܐ��s"t.~��G^/ˢ��hnh����~&ۣ�7>���hTg��(��M��N6l;���(�췿���5������o���� �����~�Q�P=�'�A���ȧ)~�q�z֬Y"ރG����U4g��gh���k��i�F������T7wK�W��C���h7+�����JCTL,�|�I���ٳG@9q�X����dS��!~|p:QT���&���>�(n��f�7����]�{U���O� ��=Ԅ�̃X{�R��*6皚i��۵ՕU�6#_�V���=C�Tu�:�(^�46����@��׿���.�����K���::v�ă�CT��6�GZ�	Q����'���'�s��[��C� k�	ύ[�g��rf|�?�{�R���?����,�RGk�loGVN��Wt�[T@�(���O���N6=�e0�������\<����l�C��<��[������,B\T8
��A^^�~�mq/���İ�(���>��01��p�0P�����8@ԸG,�����yO[�ڵk��v=^ܰ���"�Q�F��I��w
{,r���zS'QgàPU7�E�E�D�t��}=s/2T�%��9<\�4�����<��|V��ؽX�l)�������f�͛7����?�*O�b%u�Q�E����k��$����o�y��`��!�¥eЄ�l܁��]R�:{��e�u��y����4�ysfc�ĉX�n� ��[o�����4�Y1BQFm��I�֬Y�'�xBr�yԞ_�16��WFvC\�	"vc���[G��99�������ơ��$J %%�|�ь� -��c��/�)��{_ɽ7^����b)LO�Cp��˙<����ԐG�[��pn�.�c�op��u?�+;��R��A�%��_�T�O��9�6�K
%���?�Nז-[�^__/%��2È�[/��-K���1�PQQ����������B�������;��/��~�_����za�!.2f��p�NO�����X	yK��y�K���ݶ�Z��p�s�=���k����QUU%���lο^�e����[n�E�8qŃ�b�{}�gX��	6������l�A�����QZ���+"%5E��2[`Z����R<�dq��� צ�<����38�I�~v(�+[�q���ۊ:ƻ���Ĩ0vj�x^;opX<=Av��� ��w�fwbRJ�����A��]a,���a��M�J�U�g6�@9=��51ib��0�w�}����K����if%c�c�p	�����j���'��������_���a@������_5�l��48�x���+����9�v�t$%&H �5�_$���|�� ��t�xi%���>/�ɥ�(z[�ԉ)�@	[��9��e��_Cy��ٽ���k �}/r)��˚?Nb̠��[�җ������݂�da�5��?$#<<LX!���-eT]�<��4�ʚz|��m�~з�y�9��^8�zd�λ��b�hQ!8�a��`��|/=�X�D�{%��]�ES1wj2SE����el#�V}'J���T3�6a�+d��X��c�E�/˛�*\�m%Ƽ�dG��J�|qEjE�r�d���dF�]�p��ε���PX9�����wV���X89��i������Hى��N�fqb�lFGW�j�e7塚��<�Ϯ<��c�u�J�@g���>���|7?����#!2hgC����R<�X]�(Px��0<���r���F\�I�:y8o�d����g���`���@�����[�NKV#9�E��`�-=�PJ��`j��A%v�:�r<�	� .�W<�8�M\���fŹ1>�Lא�����o�i��&��A��V��e��w�8�#tDE��0�[o���n�[j��x��Mf�iSR���-�NLJ���k��yǩ�>:� uTh �Z4���`Ɗ���<K�y��w�ԩ��D����~��a㲒��v��>3M|P�r�eu e�
�����H*q��Eh������]]������J5���Պ�+gG��Iy#=6 �fD�q?]�U	8F�ێ���]|%YV*&�����h����[���/?����K�&N�uw,�ؿ|IMs�|�����������j��AZM�[[v{fg���{7��o �H�_��,�T(��v����C�!\��\�s�s,a0�w��3x�3�Yj�(R~�C��/������"|H;[��7����gz�� 3;X�_��܇c#?i��~�����m�o����H+I�3�B�:m"�v����T+�7�"W��T�Y�(��}��A2��6#5bQ���+�g�صٝ�-mM��]��ܜ�����`���5��&���ge��>����-eM=A��4{�+�D���9{&��Ӷ�4J��:<^���N;~��YAnS�pzݬ��%>�ʀ�NE�t���*��m�C�V���xlN�W��f����֣�)�u=1##�a
A[�N�?q�&�+f�5��A�/��z=Qĸ�o~c���m�OuSN��F�w˺"˟c�U����������[�m�[�Z��
u��m}�0�@�b�k_Y��)5d8y�Փ�w�=/�s��~l�R��dl$��q7�G�����M��/�&D�vI�T���Q��؊�E��	
E��A�۫�X���w2�f��3m����h$P��� H�4��e�+K�.yF�sq�6�i���kv��q5���qa�e�;m�>zW����/3tJ����UM�Uc��s����+�A�fqZ ���tKcZ� 5 |���MF���P���__�%��q��ߎK�r��o��Ʒ�\e�[@�����lS��?�    IEND�B`�PK   ��dX��) oj /   images/9b962a8e-14b5-4317-8666-1954827ef6fe.pngĻg\S��=�2�
��>zSzG�w�BT���	�����N@z��	��^H'z �����|_�{�?~��疳�.k�}�1TS]��������\IQ���z"�k����Hg����\I�O��ߟo?���I�Е���������:�� ����������ks"OOOk[W��N�<�.��(	Z"���d��x�m�{������O��݇D]kg`%��1�hU�O\dq5�Zl��|�M��l?���c�0*M���Z�ZwN��a��j�ߕ��b���������ad�~���ޒL���~0,�Ƈ�/�7d�|��b)���_N�;��3H�xg���c�AA⿏eri:��>GB��},��i;�w���J����S��E��ٮ����G#�%�ܨ�1T�{���''=���']|޹U��]�b�E�џ?*�������W 
�_@�O㩤0͌����g��A)Z,��m��ąO�s��V��I�k9y&�+����u���58����|������U�J�t�ر�����M��/���;T�1yD2���k�K�%�$Uf�U3�W$��B����K��"T?ϗTa�:�
m�p<k$��W�����YeZ��<[
�7.�����5.����/���y�_���L�܃A����d+�̿��!s��!s
�W�B.�@�r;Ku�&bt�����4��E�Y)!S�!��,�c�����aAX�J����e��[5y���F�,����f�i��x�d!H��y7��<�_�Mv�N�Q椽�Ѹ^y��-9f�q�~�q$�W�
^5?�]�?C��5(��`I�VZ��4[7��|���H��[��S�M�_�ߞ�x"+P�
*w�M�n,5�p�?��}���y{�|y��omj��M�z���4ŉu[_��'u��}�f��!f=�J/��do���{�+��鄩A��bKw��|�1e�&V�~��I<G��t�1[ˉ)$���]w�ޝ�.Γ�Y�"pi�s���O��S���ſ�2�Ϳ6��]�F����n4JF�y0lM�C��!�ު�(�AX�o�֮�Ue3#y����ٓ��2<�`�;�C2�Q��J ����N��c�u^��a�&I�^7 BN��pJ�G��i���q��	�j�tǉ�z*�?v�_� 5�[���W/���)��6mwƌ��%-[���8�.��'7r���xћ!'6^�h �����g��NS��%gvu�sώ��.��7'$���J�L��}�S�/�}ٞf��|�kb�W�)��ء杜�>v�zQ{P�uoQ=�����d�ꃀ��b����uM���պ�X*���`g���s���㍋�G�G]��H +K��,�	��RC�T(��3;��Wτf1j��D�!�%4[l�w&�e+�:��zI�^5x�2y�A�9���7N��e����-i�w���[���P�Ն'lE��)$�ɏ���S��0�a�!m�� �`D1�װ(\o�xoz力�׋��D�߁ԫ]tg�g؜!��C���t6j٤��� ���Z�=_���c#�_Q3��}C ��$����mD�$~�-��I����8 ��Y��3( �s���6q�\�1m�Rc�B���Wu4~��Ū��h��2��z�(|+�q���9�h޷�+9[]�TS�vW��e�Jr@rB�g���/[a�W�1Z��������DeL���O�OyD��u�ԁ%2�(�����{�F��lk��L6M]��8�z��T�B3�x����Ⴑ���gs׉ߙ-�^�6/�r�O�CV�3Z)�]s�P�!:�۟����C��9j��Pa�2��l��j�b���Ml�	��'9E�v7>�o��V�1���u*!�h��ίޕ��	2_G����v����X����D^��l�I�YH����z�����Yr�I����g�}Ӫ�a ��c�Nb�wO�ݝ?j<������Ĵ�ZN�]`�
(��3�i%_�F�s�� H�U\�fz��kw6��w���fË��9}��X�Rx��e�y�d'-�� ��!��;��JL}+�����S�{9<���a�0%��i��U%/�X%��T#��'���䡚��3V�[��)\f�3�H�y�Y<�c��j%��o���vR��F�4�=��K����,�ұ��؃��`�Dim�i��b��nNT�d|@yLV&T�-<��|�K�1��#�����;�W�s�^���]p�髀K�ـO��.���?��� C����kLLH�#N�g��oE��NF���|�e�����!����	�W1E�!G�%�^=;Z�f-2f
�36��.{6N�}�S�;��V�#�A��އ�E7Hx�"t�t�m?<_՟�?��D2AkMb����P�Odv�.r���c�"�x/��|m��A���f�8qr*�����b�u�����W3%^L��[8�Y!Z³kG�7k~ز
�:�S�)
�����l�c\A}�����L�׵�o�Ε��`,���|/��K�G]צ��h�����g���s�f,��4��e2r��Z~�>�Do��6�C|v�g�u뛳��tb�CeOw��]�c���/i�t�L�N��{�7+?�pя�Y�o �W�g���u����&
F�fLd��o^����>�_>�����Ċ�/��Y9dg41���w���:J�B�s��XG��+`�<�vp� �Ê��2�&����!,��nw�P���ك�-�|���n3�{�����w��|:�n�Ȟ��i�~ʑ���;�l�}6)R۹=z��EH4�_��W��'�5���.��A컬�l��_�p�}�����'����ض�Lz�VΥ�/����ƌ���+��J`�hZN¥'ŐS�f�M�ӱMz]Ig�Y�8f��]9M�Ư`�SR�`l���pA����\����u���M��#g�!H���Sy��fm������CO�-�����y��U�&��+@e�Ǐ"R�1�4��T{{����LZ��Z�ж/��}���#U���m����:՞��g��ɫT��k&N�詝O�#z��"{!�زw2�n�r��<8�c�]jǼU6�r��r�>�J@n�W*�U,��|�i	a����˼��oB��~|I�X6�h*k:���݆�Q�G�M��P4d�3s[p�Uk���qc���X��ں���cCs�J�x�-R��tojg:wt��f|�9=�c�a��s��J~�RWs���E{"U�G�����t��tj�*��
��1ũ)��1M���ԫ.=��T�㙫�
����q���H�-u�H�0=¹@ؿW�Y1��JK�:�"��J�\=LJ*',=�g�G_{���I�~l�b��w��G�\��Vk��=�juڡq~�˪��:w�q.��&*XUz�"�Ķ����ι~}kI
�w�2�^��>5u��?5}��%N�*�@R��}1x ���4C+�c�����i�Խ��*/��3����O/܆�7�[_��W�).~b���������72�}_0������-Zluq(���*�Cb(!���G��.8[�~��ɑ'�y�#�N)Sh0��wЦ>��� 9�` 4%�	�m8+������� ��W(��Mlg��f�z��D*�-�ӗ������>t�5t�IO�]�v_w��DA74K��u���^m�1��q�6��xp�'q=%����AP^ݘ�ݸ�nt�t���t7e�Y����^r�]n�b�f��[�¡9�o
����8^հć#n�w4��*�}n(���r���Q��U���i�����8}k㟜o�ש�>y��,�;Ѧ��b�y��]z)�����Zo��n[g4�zٚ��ܖ��i.��[8��L��1�r
&p��{��2���/���k��G�I��%0R�ۘ]� f
�}jY����9�a%�2��]�0�Q�������k|�L��&�Txlʹ>��t�&[Y�ar�}˰�����F��q���L&������;���/WdГ��Z&��N��|�d(j��-b�r�^Cֳ����ܖq��V���|҉u�:>Hf*��e��벤�YZ�3BS�����|JQ��!�6;^G�#�g	>�v����L��yºL_�,N&"�����u�Q����V@�w! �������m�*1�S*,N1�g36�B��J�=2�o����/�
��L��}H�����\��+���������"NwC���-@*�+a���&�({� �����x\!���ԖJfc�ݧ"lL�J�R4ob�.��}���I�d���d{�DB\�l[A.�k�@����0� u�D�	��y�	��	w��[��^'�r���	�ƎިC���Y��B������/���P|��t��y�d��Y���)^6�{�:v@��t$��|�-�&.r��>� �L�zGjv}�	���OgFq��?6jF���)�
��::ߝ�^*���Fz��nOn^�8��W.ǭԂ��0L�:Q�7�<�~���7���t���эh�I��?�@E�?�o���v(:�����5���󼳈UW��P��Ʃ�8��~��h��YN�r�Mi��BNW\D�m}�θ��a�c���������}�)z�l�j���-��1S�;ǣ���л-�`"���$�.�x)xi׵!�rf�:ޗ�vhVLdc2# ������qiݵn��C����7"s�#�Y������lR�+�0)�Cݷj�yK��I���TgҮ�䮇'�a�׭=Z��ўL;⸕*�����@�ƛ�~���-�-&JL�ĺ1�bC�D�r�0�%��~�g\�3���=0�o���=}JEE�ǃ�3����'�/�p""mO�6K��((;;���ar�瓼�B�r���^k�����7���?�\&FIg	|�958*��Jζ̩�GV��!��8�v7�i�P��jɯ��z��p��7}/E�A�W�y����ѭ��D8e�S���1�]t�|v��w�v.`/�Un��;�U�P����2�d�����;tH\R�4l-=l��dZ��(��{��^�-��2��(���0��0��CF���������J�--���޷�_h�M��I�ޭ���y\ ��p�*a�;z�K�G���?S�B@&r��RC˟���v�Z�$�\v^��I�܈n�;[��W'n�~�@7�> �b��4�Kdq��[�2|t����蹃^��6�JRp��@XES#���?G��:�{�*/le�W����yI�u�	�~���VXכ��
����~Үk���['���1_3kO(h��4�Wۍ�$�ac�|�>e�  Ks�����'�c�6w$_p�1���c(�����~Y�u~��i)lG��k��&w��',���B#�ё������m�u��D�!)�]� �>�Z�2�>�fM��-���d+���v�����+��(��S6�X�B����"zLycC�рLm����7�U��0_��l���~hH3��N��JD��1aP���}[z�W�^x�Rt�;��<g��2kS�V�g���W�yꞶ4v�;�\'��w?e�۱�]C��{S���17�Q�L�����	�Ļ�y��\I�y7F�)�uk����X�D7׀K��
�yQ
��ρ��rXpm[[����$|<{�ߟ��:�S- ������� Pe�'|�uF�*:�"�6��h��6��w����:��=1m�ß����-��"7AՕ���Q��/��s���ve+�/JԣM`|��f'��@����� -��͎̀����!�w���'�$�>@:= ����F�Syy�3��D�\	���C�ʒ3�� ?_�U#���g]�L�2��n�~+}��ח8_�o��a*�X5nSD�w��s���g�"��~�i��ްO�mLs���l��}�WyV=�^���(�*��c�Yy� g��'l�Cl�M��X>�U�.�\C��+B���hi	��v����{:&&�[ȭ8UsC�@�L)�P�6VV�<��Bm��y��JߑXXі�`x^Ͳ�Ӑ�~���x5Ke�޳;�F�	"��k�BGJ�,�\� ]���b.�aC�ً.��s�0��r{_��8[� P\ķ���������ʠ��+���f��k�a�ݦ��!Q�⏐
�pAMދr��k�&��%3J�7~�%��f�n���ښ��.HI�U�@`3�[���޷~���9Z������{=��۾�i�9�s����k=<�7���8����;�!�~����\g �D�筕����~^ѧ��{��"�H)l��h��O4~|�n��?��d��a��HU]�A���L�k[�]���_g5&�V�q_�|��S>g뭿��a����U�����9
���vp={��O7���u�ѯrarّ��ѓ��2[%Zmk��_O�l6-2YTD�f�W����g�+�q�w5�~8���8�nD]�V�Gv�3"9�,�M1ar}��m��E����"�{Y���Q����6�U��U�,ܒ�#���t\�dU7�`f��ҫŴ����0Om�e�:77��OC����$W��=����x��{ �X[~�2�f%�8xO�X�[��-ADV9o��D��%#�G�\�3�LR\V�c�N��}������Ís�RuY�\;2Tb�ǚ)��3��V���I��
Q��'���5���F�&
��$'8�f���A��ɄD�ۑs�I'��𻛺ƵVJ�M�?��U��Ǜ'�1Hp�<�Rݠ�U=b_d���)�Rf_�L%|�`�=�]���,�+��G��&��F;5�,�Z�I_X+q�Ln��ޙ�~�|����vT�5�S���v:�P@皂�V�>ݞI,Iٔ�"��%塡ɬXNgh5�w:]ۢ��A��*�*����Z@����H�L�;Jt� ;[ ��4m���N��6y�U���kq���7��������8��3�m?l��'ޞ���j4���g���b��s�U���97�|���`�{���2�1��]L���)�6��k,��Ї�:å�ۂ�<U\*�55F@�3Y�_\T�g DD�a���ɋ�����\^N�.	���^0�^�R�����L�c��9��S��I��}R��ӭ����iX+���~�n��˵�
�/c5pgS�r���9���e2��!�=�#��W��j������r�]|��>Y7�\V����ɪ����[��m�J����u� �r��@�1�6�1�ĦX�<��`�e,2!~d���ex�b��`�ܨu.�{�h	�2�9NN?�'�S^B���wGa���3�9��ɺ��PBo�9�ae�Z�^8�(�``��e� m央�Q�G�T�a��� ܌���Gg]0���^!���k�+�U>�kvWx���l)��&�X>��j��7��e&�<aw L������>��!���S��B�m��G��>!]��ʟ�j�o/�PQxQC
e�/`jS	?;l,07P�5��a�ѽ4���o��#P��bwȂ?[�l�q7P��'H��G@���_nشS�FR�ZJ�[v�vO��q:@��u4��8�3�4�z�f�����\[S��\YCW���0T4z�-�U��J.G�m`
m<����e~LoN4 1�����5��j�pj��#j��x9w�C#SA�����
K-�xN�.�K�i4�o��(��D��٣���K �dP��Ј��{6��@���lʞË�7K��*����@������'������:�*�mp��^���L���Td���
�u� �n{�f�j��)�;�d�4��Ƚ��6MQ4�
AO �|��\ݸ����lD��ig���o���Tk�&�S�q�ǌa_�p��Õ�\����d��aR$�buچ��]q	,ݏ��4�6�5އ555��&`�@��8>�.� ��>�N鮸i���Y2�iP����c��<���p�l��;��&Ӗ��=�	�EB�C+no��Y�ۓ�<����J���*�l��_P�P$j2&Vr62C�ѱ�m�Ĵ�d�ׯmn�~��Ͼd�Y��I�w���H����ۃ�z	ey
�xYH�5AIM�<\�J�Bi�9����SO2���J���u(���U�fC����4�]V�o��������J\xL��j���o��wg���G���tL%A�X
 ��f�-�]E%wa��lq��9�ҿ[���c�]�� 8���I(5��b}c�4����/;8덧�G�џj �~+�6��?�ߜ�,]8�Ձ������U�MTd��;F �$v/?��&t�z\�2@`q�|�?�g�.����Ϸ�Y���j&�%����yԣ�j����F�Zw��C�������c�-[
+�B�aUE�S�<~j!m¦�Wb���j�уy�K�vΎQB�_2���H�`�|mh�:�^���zA�Զ���f��Q4������|���<Wj�o#���zNm&��	ͭۻ�k�����o�x�=��N�pz:9�9Jh5�=����&H��z\�����X��1��������s�S�rkF�	K4?��c����]ߜ��˝��v\���ޙ7s�\���#
I��SSu/�7V37�f��ǣ	���	�U,|'Y��8kd?W����������+ ��6"�]o:<�]�6E���+류�I�q@h���Y���{(U-�ʤ�ؗ�.��R�C��q�s�e���"�xr��/�<X��.VΞ�6�����|����%�\
Ҿ	� ��O�����Te�X��9��%��x��녔n�i[�)���El��4�����[��u��ae
�SVSX9��<�Ǉ��,��	{n48$��K�T�G.�D{{�k�����k�mG;��F��|��2i�m��r!��N��2����.��?-�a�C�s�,�d9��y���G�r��6ڼ�>:w�:�	`��H�Y����l��#��zxdZn�Ď�y��X�:/��&���%��0��<X����RW����s�yK���L[Q��/�ϛ4�6�-_�4W��蓡B�>�ΰ��۬��O�QI7v��fKh$�be�����ٺp��z�����WA�)�����vH�h'������2�bz8�F�Y\
���wv�j+ʗ��LM��K�<d��l	�j��ى��C���&�W52�"�J"B�'�*-(��tR�����р�L���5�"�~�'UjZ��j1|9o��dT�T� F���P��`���.��e^O��Lk���w^;�>�*�=�b�����+Qn�N����Z����&#_��oV/��۩���νKZWrB�A ���w�b��I8{=I2�Bh�MM+��vu���8A�ˉ{�δƓ��!I��풴| e��U�{��Z�£+��@��o��B< ���H���K�s+��R/pn�@�-��cִ��\W:�W�x����=��e�1�g��Y1~���e�$'=~����L|�d�|�~�/����/��̘V[�kmCKe���r}s��_ӥi���+�م�Z2H����v�ϒf���g���b�V��0���H���ݠ�H`R�`9���ۏM�o�z���,U��%G\Jt[�:�Ӧѣ�e5�0�{�Oj����7OJw�u��8}D�X��(?�d&���{���`.ğ>�;��Q}�f3ͣ���&.)��#����+5.�J�A=�o��o&��,V���Uߘ��5*5i�`%��v��z�;Y���C�Nf�D��{�SV9w.u�������ĝ�����f>B���^��c�����!�n���O�*��%8�UO�������S�'��6H�,uO��rG��.]�t*����a�_8����ky��j�琎�
��7�\���/����_*� �o\ҥϊ�s���xr���!U���0��������,�`�.(���A8��H��B��*<����]2v���f�R���t����*�
wqO�F\H_��I��R�;W&�g�	Cq�,|���U&�f�=�"�݁��W13(�����=����!*�z�h�I����Cac�Ϋ�m�C��3	�Y{��@]���u���������LWZ���p��Yc��;��|@l����*�/�*VC�v��[��)Z�`�ӝ]��y���׏�ofl��e5��d)����PJ2���󰜙0���Y�Mݳ0��YQ���㟀�^b���|j888X�ZJ��&s���x�P��b!f&w��a�`��	v���}��](�q��<Sx��t�-��
��*�QU˲�]��ˊ����W@��dq�]ۇ�������N��T��ap����4a{$#��ʵ��#�XP�<$���#\@�8�-o=eT
���Ĳ�C��FNx+�+֓}�)&�M��/���8�ш+�X�����!$j�=��{�G^�_ NN�~{5���R| Zvg��	��Q�3�h.X=Lf���ߌ����lQ�=��O��ٚ�/o=���ӳY��,	�g���s���3�M;S3�*�9bS�i�>�OH����3S�Q��R%�vdw�1PX�.����oD�D���a�,�g��l��U��IF����5 ��}N�!�R�V��Չ%��c�$Se���Xy��i�}B颋m.��� d�2U�m���#�)s%�}���ˏ�O=�u~�z����=�81�$�1F�P̳267�3Se��1�,����0��'����䖅����D|�(�l�?�f6�1�����>(p�.����1E$G�<A���p$���t�����w���QNr�nAY��s�I�Q�)A���������F��i��q�H�\+�wi%9n�'qU��%_:�d鍋;W�c�?�q�5Y����k���c	۷����t5ޜ�s ����H��bH���Ÿ�.���Ƈ2�x=��zV$!�{C�r�y�� \��<��{c�_dT���	°�ժ;�py��顺��.)��םO��b̊�V�Yn�Z��0Wre#b$N�k6-�+3��?��%�*��d�!8UH]�w���z�ґ�Q�L�a��$�T�A}����E�\ �Xx����?C؁����bM@:�}����͚<�/����`d,W��(��^:�s�	i�V7�1e�\�c�l��G�
�˰𓾰&��{Ҁ�q����^�48}:���j�=���X���3�ڴ޳����:l[���w�o-]�����i�-T7f�{�t��~�M@g�L���ä������+���(�u�fվ��2[^օ���{d�Y"�0����I����!(��P���|�IҠ	���R���o�~�Q��,�4~a�c5
R$�;�{������Mռ�u�����Z5G�xE�������a�/�?W�UIy�#����@]Vb�����B�OK� �/�����6�ɺ��<x�d�@ �Q��k
�Nv.��6�Ȇ�r��t�۽؆��u�*6�YU�_fk��������C����Q+����6�ɾH��6=��Ǿ���'3rvWk��x��O�.���{,��{�G%��C{.���VF����{� :��_ʨ�J�#oPo0���[��HY\��i|(d��+��8��D'�PKk�Gٍ�jl0����2�ڱ���a�C��Z�km���&�}Z�?��v2�>���߼
~��5��g�;�#P��M	+�1���9��z$?"����΃�M��/��4�{�*.�Ѐ�����>�S���W��I�wy�r���y�^�M�K2 �NP�q��!�Th��͟X);��ʗ�H�`�<ᐾ�[�i��'f^�#�R}z�(���/kE��)7��$��ׅ<��[)�
�֍CJ֖��'��5�3�j�lPs��K��V��aO���l��YO�|��O|r�5Ua; �H�-z�a&�W�sH1�	+�#&~A)�m+�vD�%�U}��z�mN�u)�z}�l��
K=o��_�_�?�OX|��ǋ�`��ir��$�c�]���_����k#��h'���	�eS�e���nB���4�&#1Vۍ˶��I��p��ں4GIC�kc���C��c��8'��b���`k���������F���.!��N�vM�r��v�\>�Ą�7��M���w�Y�f��v}��Sb�'V���͒xp�!�2xUU����a�~V����gxX�.5�S�?����r�5~)��֪%�]{�+鼘�7Ӽ?�Z����G)iTOb������������(.Y��ŋ���P��dڬ�n��{-�	cݜ3��Z��3�:r��S��G��2#W��
��jk9nF�Qc9��lR�]�����[{Ψ�z�?���]4|p2��`EMbI5�B�+7u��fɝWР&'iֳ�7���bl�����<L�E\#h^=��B�����_��;���^Y�)`��6d����֕^����r-*�j�)��p����ϔfH}=uH-����2Ϲ�$&�Y�x}��\j�F�c?ơw�qP��nq��/���P�fs]��.����ݞ�q῁Qӿ�;'�&t���o��y���6���|��X�p�1C�އ�K���9mK�����P=���}_/�� �u(�8/ƼmNV���t�D��d�ed2M�k�0���O�N�)�ք� �ɫ�k���Q���M���js	�vU��7��b��4Ԟ���#
�Gt�B]��o�0OOx���M{_�3tw_��w�`�>v��/w�it���J�N?�2���	�Zi|�:FR�����7`Z`��?���*�Zn��F��~a����{8�X����=]��#zh>�����Ԋ���b�Yj�#�����g
.�RQkB?.����|���]p�g<�����֓�׬_	T������2b!C�E���x	�^�U��/���m�j22gՕE�����]�B?�B%��J�$�j�����,�`���}�4����<ӎ�Z���&O�k*TՈI�] ��Ӟֵ�/XA�=�[�`VN��f�"<���S���ه��b�w��`2��.�X�7�Rm�V͑�Qn����V��x�G�������o����z���|��I�?�(�ܙ��¯t��OΟ/h�ǻmZ�.���j���?���*�%�ʟ�4L�.#���RVE�s)77Y�s9����? �io���X��%�-���x;q�p�ˣA�ҋ��v)?
)᧻����Z6V0��\��;k�( �x* ;NvT��_?=��^3�xЋ�*
 (��(��m0��V�1���)�G�;�Տ<���t��'�m�����a]�|�hq^�N�	8%���Q��Ur�SF�=J1�p���H�0��m���o[5sg[�0������_���^�뽿�_RV��u��	?D��U\���_i���N�0�v3�o� ��~�ɼ�
AR�;�]�n��?���
S�N�\�
�vt.P���+K��?�_�xnb��,ȹ���b�;y��f�����Uǀ7��.���(����HQ����ôh#>b��u]L��a�/��fx��"��L��<��i�!N�e���X��2>� ��V:��3v��QB<���������A��z����!!o�X�\��_hPIE��Ѐ0��}��Gf^}��%��~�W}D�v��t����#vy�Rh�?_e�*�Uv�8Πƞⵝ&1S�6��D���n�$��F2�׳�Gقz:q9��k�3�:�}9Φ��>fmL�M@�V8̏_*U���?�;�nK^��y�-֤�-�:	h>,�w�K�Z ���}iwǡ4Q
u�K���%�"j&��t��O
�6�����v=�8���]\S�HŔ��[xzڂ��[ג�H�$?�Hz+��$����÷�}yt���WC����ؾf�^E�+��Ÿ�j��d���i�]�I/j:>�H�����3�B�a?���ۇ/z�k�:M����N}'���6�<�M{�H���x���.;B/�r"��l������O�c�/�H5OqzJ;�|�bSN��#��0ʺ����z}3�6Y��y���\��:�L�Ld�O__j\W����"WWwwrt�"��3�B�����_V���bV�Rb�Ѽ����)����az,[]`���s�}��$>~E�R�=��=3�޴���/~V��e�g�F>��]��'�MM���Y�|����^ѧ�Yeoʸ:iA}l�OO���~�uB�9_�ڊ
�r����I����ݐ�<��'�w�n��?���=�}�U���EH�%^�D�4-L��NS�%�Dg�T~��6���b��rl�ê1]����R�5/G�#�O���B��vy/��K���ϓ�|+���S65m�!�37�S���S�,�3z�
4p�Q�]��!�o���1��-n�IW)�g��'�|���'������{<��W�U'���K�1���k���kc By���� ���KW��ge[ճW����=�WQ�e�M����Ǽ'�Q��S�����mUe���@�+��ѭл俆�㲲�߸qC�g�q�h��o�ݏ�%��Q}.�T{�
�6�R��|�yk#1#����c�W����.f���Qr~�����}w;�n��\$���=�*��`�2���C�-��x�:)OjiTd�"�>,�}�_H�����p��|�������~V8o�6�^�u��ߵ9�~�
m�=�Xn�Pm��q2xp��h�霺�t�-��}_�}<;"�W��$�bl�q��-�E�dcs�rb`\�󮔺����8���^B�f�.�Ul�,�>�����{���\�ԛ���U�%=Î�`w�zGH��=����8\�2�?cgz�Nã�tx���_i(��ݩ��g�S�� �τ�+�;���P�	n]�ҧ_��6N�9a)!�mu���k��{ɾQK���ڗȑ��DP���#��I�^��b���T�{�Q��[ʥΟK�d��	�h�?���5T{,L	�N�GG~�brS�\��w�xyҼ�_�����F�u��4~�	W�A>�����R)�_ZM|Y���x��D��4��C���N�>�S�ӛ���.���wo'�<[��|֥]��ǁ���<M=�[)�ܙ��.4`L|�N���U��-�Z�Bҹ:{�TGa|�e��������vά�])�:]r�p��3.3�3u=>� ��{_,0����&fͻ˞��&%�/�����!��������D��o��a���)���q���j4����	���l�u�$fZ�_�+���eRW�|�������0�����sc	��Gb&g�q��3�t�򛿼�Wi�7�E�b��$��;���r�U�b��{�*Skrپ\�m��i�u�.'>�0�b	����',>�0�E6�|W���6�P��#�[�%4�O����yX�����2>k�D�<�����uўs�
?�.��-�����t>x�h��rҴ��a�f�)HY�o���;�
ϑx"U�^Ys�H�;�-����C�<Ðk�B\VKF�Ya�]j�u��t+��H1|��i�<v$�]4��S��U�P�9WH�?sn������5�_����bO��~�n�r��jF?�_p�`ۈ0i,w���`[%�����������r�vڤ��y7F.�Ky�N?��c;�^��D����<�� �k�t��}gZ|
���vv�8����߅"���N�_�^��b4j.42��c7h��CL5��K;�ɣ8�w?�u;btK}*��O)\цBu�c��cz�o*N\�ku�������3��F4�?)���ԇM�f�D��O润��')>ʴ�x{5���뫍W�4��nL?�tq��#�6�i�xy���49�}pP��^�+f?]#u\���s��a�1R��'����x�~ay",�e��g̶�'���;[�S��{Mo�ɀ�df'���C�\ӆ}J7�����Ơ){��[߲l)4�s��'��)��UA��ύ@��JAb
����b�
2�ѓ����q�:oi^��y%���q�V���3�Xv�n�^��_��-�1�!���͸��^�P���e��V����n)(�r��w�k]|t�mdP��>/X74B[;ܾ���	@� z�z.Df�}݁Q���n��IA�Lg;�����0܀�9�w�W�X��%#jv������C�aS\�f�������hi(ɯ�Q�5��6$)4�|~��su}r����Z���<r������י-g��F��_B;v20�ߚlK��E
>.�wS��?}�,� :0Z�}4�� �\��)>�o������q�㤥U���<�fX��¨�K��[r��S꘥�ƶ+-��1:�s}����h�(>����1��P'��wa�s�����q-�JӍ��uy�t8���$HX��x�P�o�7�k�U*��t)5�o=�#���Uǘ{������^dOB`n�����3\�� �ڶ�uZ�v������9���c���w��Mn�
�J͸����]܆
��^��7��L���]�f���n���C�[��
���!K�����C�y�|]|�������ѩ�z�5�.�ů5]̆w�)��[�xa��&i�[=����vW��[�ǔ)�{�LX�������\��M{�_�=�sx����F����5��!��]�ݤ�>S~�K^��u3r69��5ɫ6�E=����mv�[r��V+#1_#7�����J�1�,�UFD�ȳ8�ͨgs���=&&�}|�9�w;�Ь�ƽ�A��hR�K-�n���E����,���Em��e͘O�>P����{�Ze��?���q�<���(���f�q0�KV��Q2�����]1'3��K24������$�*6�c"V��\�SέkG�-wwhQӒ�����xX4�,��V���Ӎ��Am^��D���_yVj����}��O[,��1%�@q��Ɩ�Aa��Q_�����y�;~�_,
/�(8�|@`7L��PW��@��;&w��^t#���,��<(��h(G?4y
�7����Lb�I��S�7��(�_+Z���F�0\�ch���z�xc�=���k�$���k�����&�A�CB���A������S	��;�����Y�ߢ���;���0�����\׉*�ݒ��ް⛹6gv���5D�bO�!OҜB�߯�ԐT�B�\߽�l�ȢW�[�Q8���Zk].�p� ���\"�G|Q>~��s���C���Ć.�tD��;����.t����\|������d%N2��4����WxG��]�7B�_���4~���ax���!��BZF�}U#����wϊ7ڊ��s��wM��[NԵ(ԤiT_��4�$���Cr;����b�W�������B���?m�/�{��'Pܕ6��~e�H��{�۟_��L�Gpۂ�Z[��z�YD µz�hT㲷]���b�v�Ma�T�M�9���C��C�@��c��J�KY��yH��x��-�h�\����˒��m�8�r&����~�ގ�j�G�*�d�qB��'^޺�M�X�y�f�Jg���-y�l��5��_���UxU��9M<�	�f��c�4���I�V�!V����`��"�B>ka�-������%LȬ�h�S`b51ӥ�y�7;�FZ\�
�#.�S��Q2�� Y�k�>���@�E�����__���}.���Z��{+�:��
!W���͙�(�r�Z�0�^J�����/\[P��h�lR?M�
ZB䑬9��8Y�ۚ��w}��E>�3����x�8�81��wQnn�i䷱u�����z޵�3�Bp�Z\��e�RP�0�tw���8�y�t���K����7 G����x����)�p��B�q� g�;������������Rg��7�w*�]��!���?��E	_��t���j|R���	��q^�6o��SΘm�5��r�(<M`�o�s�r�!�9&6��N����+�{Ƃ��K��N��Y��5�CfL��Θ�G������b��&��]������qO6��GƧ����e���U�ϕX\��>R���p�NW$M��T������>���ړ��L��@؅�d$���Δ�Ҥ:W\Y�4��m�v�|`�[�l�is��)��*�^�����+x���%<%g��{����D	v����Y��5!���Vk|>��c�?�q�J�I�q쩕�㶉%���������^�*a5h֨}u��)k�yc����0kv������ <�$-8�~��پ�9ލ@or�8�fCH*�l�]������`���1+L�xk��M��u�o����.����?���8��w��m��*.�k��	��[*�*R�������v���bv�Lm\�v�	��熥����wϖ�ֽ�gZ-�M&x��*�̹�9m�e�.Q��$��l4�Up<v�f�4ġ�"_F���-�)v֑2�C���/,��0�������zRy�ɩh�6'\5�U�V����IV��!��@�����l����Y$+��`�ݪ���{�(M��Ϙw�wk��ri
��~��K�����\���T�����v�cf����e`��D�\�5�I��z�������8�{�co,E]�<��o����S�X��]_%�_���$����D��f���̂�L�` ��?��з�����S\�d��n���ߛ� Y����*6h@/�{m�-!J��~�
5l����g�m��ւ�c�7��[|&���ה�isC^I���f���}�#�hHVr�1w��zgf�(Y����5uUf����K���q�K����u7n"�V��}y�y�}!�'��������4��p-wخq7ܬ�S��&އ]�UP�~
I���x�jC3�z'��y"9&�Lb��e�V]�]�

���$(l]Pm�ē*t����sw�ur���(+W���M��*|.KMQL�@H�ztw7R��j���mӹ��Uƹ+�K�|t
@��t ;��,'� �n��2ŬKZ�kL�=��th�L��\嶕tt������%[�������VnR,�'�q�)�̟���u(���b�/�����sr�U_K�(��~3*1�z�v��l��c�s����o�|6)�~a<�Z�F¤������0����Q��3����鷙ߪ�1�(���A~��B>�"�~2�[.onU���;~\ƭ���u�Ga��l)d8��ψ�I�Pۖt���\�3;����r���vb8m�7*����Bzi�>�4�Ĺ	�65����hZ�AZ�ڑ�#����ר��n�KJQ���/ú�1O�'F���!������ �781,��.y���F��:S�"(����8>�����''��-��3��Jv"	�k�ר�֗6�.Y�7�>/E�N�Cg�&��9)M�h����L��[e5���q����?�F! �<�g��c⡸c;>Nd|�:R��x��"�+Y
�	kƬ!�����k��n�޵����-�?�;�@�ԭ��k3�x�ѻ>��u����b"Ԩ?��q�3H:rݷ�upq��È�����x���u�`{��`���q�:���he��+�Ն�,u��c5�,��US*�Ō�=�r�0��L���љ�N�֮��/�o�"����� ^f�]�q�-f�tl���5�� CM��M�NET�Q��T|#c���@FN�|4�O7��QDDDp��gL���=��gޛ�I�ȵ"7a������%aI��2��O6���gغ����a;�U�9���Q̏If̋��|���n#�}�Fϰ�%W]��m,U\���׿�������mV@O[��é���g�����D��D�wEBӿ�/�`��A�G������K8PgS�(�}��)��..�Ws�^������[��s*��q.[�����	����ݮ�b�cB��Ҋ	�>6����]ە$���N�[�Ǽqm4�#0�S��Y�ed�44�rhY���*�"2;���	�Ф������Cea�}�aRO��a�0�F��:X?�s��R�?i^�9�����@
,{$�z������S��rDiހ(�D���50w����N%�hE2@g��2Эwa�!�n�wΟ/	eu�ܹ��_��O�+�cBvU���/��1ש�_�;�� ��<d���/����g�V���Xr���&���У�������M	�6D���.��ll0��C{�?竭b҅���G��-7:�4�?u����S�ɷ����HQ� ʄx�|Z&u$EY�TN}ϰ�CRB��]̬�ٵ|�&lw�vK�S�6�k�zʁ�r��1vG��eҘ!T��ӑ�ɞ3����Q=��!B�nZ��vZ~bL�ro�q�v]]]$����3���M^%��{X��v�������)���k���}/��z�G�Z�4fu�p���72�]��/ ��'�Xu#3�P�)/q7�6�"k*E5��/p���Gb���9�y'~IE}���:X���ڨ����;��X�W��f�p�ՙ{~rZIӷU�j��)�J51�;mo\o��R2�Y�{�xR�V�����d�YWiQ��vZ���F�]頃�UB)��ue�m���!ϚC!X9Z��3c�y�?;�r��;4���o�gN��ܔ2�T��?63���-uBu�����*��mG�����r���
��e6��)ϑٴ����ǂ�F����|���]8��%`K�%��ђ[�O�V���^'���8���w �J��Ȧ��3*��@�S������RD���� �˒6+u�����T@�%2�YC4\M��񢢖IJ��C��\��e5a��,q��]�{f������&=�����*\�/�1y������Nx�sVjZ�:2a"����A��ba���|����� � ��UQYp����r�������S���[�.2b1��;e�M��{q��z=ߟ�a�l��*��^^���׶Kx9Ԉ���W����$�������������KҶ���M+�����.��p:�&\o��e�?�����|1�?���A�|��(�ZP[��P#hځ�c_���ٌ���ռ��a+���ֲ�?��!<ɋU����D����Ђ��p˛����kt�a�ㆵʤ��R�,��H�	��Z��8����g)�)���JOx�P���n1��ف&�$)Vof6��+�A܎�?��|�P�2���ԋ+�n�Kˊ�^��/�_�j�}�S!'P!�Xϟp)�tw�Q��Cx�S�d�j$��i���㝺�h��N��� �Y������ۏ�m,�a.=��N<�XЌ0�54�}����{�L6�І�Q�^_M�\Z׿$|��;}��N�0C��,^͋�k�C zgW���5�)�j���fl-$Z3y�(tFT��k���!�h�2&{�9-2�����1'C�CE��u�|��gE��x2	"�J)���u��Ξ��;C�Y��{'|l={�,�������%7�Q�c#˽F�9cw���kɅR��/��!Rsoǹ�/�&ٳ��!\��X�#��f,z�s���/�Y���6�5u/:�[4�,�����E��-�.��d��e�J[�ߓ��܂^b��O������:y:���O�OgU�#���f���4��"�݂�|�|�7Vi���w.`6!߫�rl�m��賬�{�bI��"sB�y�hȆ$�?�����"(�޼TBA]`�X��/���,b�	=�:iq5���c��hږ I���y^� ��)�}�^���?���L^��zv0�z�DN�<{9vv��Y���u�aP�ƀ���tdѝ�1��ތ5�(\��?�h�C3g�sM�$��C?a���
��|��hG����{߿
���������w�w�fo7�<�U��d=~�r�V6�i�� �V�c�j�^#�#�C�
�ʑeJ2�r&����n���1�'`��z,]��A�a���5ݜs^U-|_�G��b�p��y)��l�4�&�B2�iQ����9}!pS���O��=�Q���Xn�D��,��o�z�[�]TRs>����z��/U�����+ދ�>�������ן�8�ޙIƸPK,�3P�#�1�m�i��=?�H���"�lXC�O��R�x��8�����v�_���<���:<I-��2J��^e�(�O:a��;$8�:�p�:h�+��<o�C:f�,���:W��;a�t]I#���A��{C�/��й\mnY"��0w[: ?�s}�9�,����.J/	����%����ӵ0\��WN״��ǿ�^q�6;D��Y���/�9����>q�R�����y�UJl9[���R�B�L��X�~%o�Pgi�t���;{Є	�O%nud�ʲdn��6iC'�c/��n��g�&^}_������8�/&���(X�����2�H�Ȼ\�O)����y�1y�|���C"��eq�L�5S�������.�����?yx�Qq���h��d�Ui6p]N�mQd��o_1z����+�vYJ�0�u�[�i����6<)���G�2v���� ��`2O�ڃ���bÎW� �F�y��&�t��DP��c��Q~2�rDkb�͞^gy�Г4Ѝ�*���'�[�"�����G�����@=���܌��D��6uT�����z�v��W�>��_�$���IY�_�~�P���>`�u�p\����&�v����%ܶÇw .�|̃9�~�cBw��U6|�,�a��ئXWx�f���(��>݄�gOl�c�wO����ݮ�&QaEY�l�!��k��?[u+O�A����Vv���%C��Y���'���1AA���^$%{�W`���sR� 6���hpm���H�m:����j�-�j��?���dz�;�#��|�j��ZAp�!�FB���z��3�
�
ae��fUb�z9�b������S�cd!ۛ`���<�v��=��g�#�.�n�f[�OΙ7u�G�f�.��#x��=��������&�*�+ⴠa�opa�,Kp�E��m��ߴr<��8r r�SY�\��tn�����7��v�@���~�_�4�����֊<���3̒��WPN��'1c4
1��TҎP�Vf�]��o�'-;�gw�p�с��|��_�nY�}0~hRme����ѴHڢ�4� �ǭ0~{H��/�|1a�X/��(��T�I�s � �
1?�k=04i@����]~ƚ�n�,y۾/t�V�f6�.<��_a������-�z2��5���SI�Zx�z���L%�0Zx��%��F<���;��9���� ĩq��J=P:K�$�|V�b��z�6v}%�ni���X '�~Bp�.��'{��e.ᡝ��{|���e��e)3�x��SY����HWb�u^*��|mJ/��ǣ빅�53T��cc"�Y�RQ�!�0��t�!�-��<b�"�]0��_.�9��^�֯'��$c�^�u$��)l?�IN�5�?��.M�S-��ȣ7��Y�H(��9�01���M��:	�c�����%��Ҙ�h������a=� �[��߽l}%f�(kF�q��P�hq��f{. �M��d��"|- �/�k���-Ccq����(h���W�A����`(Pvu-B�a�k�Hxۻx 	_��+<2B��ٿХ���"G,������>��n�k�ׄ�*�ί�0���U�0�dwz�BH�?�-j#��rr���/�C���}�&{�㵡c;hB�	��tȣ���0a���\f�L�܎�Ƈf�A:�=;=3�������>�4�9�.fgl"�f�x��賛o�ۙ�F�~��-J��F�>�6	���T�����B�4n<$�_=+YF��\GxN�L����pUPЁ����p�����>~�8|�j�,L���~�^aS4YƆ�����'�֡�Dg��3�WHX�^����Y3�[n��1�"n#+�Z��׎��H�(��d�dYfb��2	��&��u���Ls�i��1)Vzd�2�s��d��/�>͸ل���r�0��z�������������F�9�5P�~ʟ%&��{р�{�Ӣ�˥}��~�4�u�8tI�U$����~�m+�-�� òh�/�<.1)���JT���L�P��|gRAv����m���"�m:x.l�B$b4:��t��x^�K�	q��]>�Z颎�/w�g����̩U)���Ƨ#�U�17R��Loj��/mz��YG�������\/�N.����ӻ۝����K������zOd������￉�%�M}�Q�p�O/�k�����A��u�6o�g����~T�a�N�VI�b��"�Od;�Ϯ� �w�A�G��d�����/��ߠ�F2IA{��V�2�n���jtzU�{8*�2������iK�%J}���{2�{g�#�@u܋�/�'���)s���d-����.����V�д�����ZM�9!<:P��t�>=�w'����A��P�� �D����R���d�k�
��31�ܸ7�"c�/�G��TbĬ*m^�R�}y^��LL��f�'K�И�94�P��"�\��j�O�_�>��a��tbJƄ� ��Ij7�t��@�ko;�pZ٢�6�*56$�����*�U5�|�O�o���5��m\���<��s�5��n�?2�Ni����EG��h}�|�����3�)A�/Q���Ң>���6 �l�tx�1$�}������c��IsL&H�A�"Hj��5�7&��o7J;.��;q���M�2ǧ��{�USB��'�O�)� �L�Љs�ۓ7�I�����d=�.�d�����5�c����ِc��c�7�8�Kē8�\}�����s�ګdA5`���8�c?���>�cxJ�s�6��e"�_�$��ޕ����Q�Z
8u��Z�'-��J�#z{%S*�0����M���ӕ�/�6�4wuf�툦s@)I��/�{�	�)�z2�S�j�^��d��\~��A: ��$ʺ��׹��tX���l ~�]��\�}F� �ǚt��6�;�V�xED��8%��g(�Y�Puul�S�������&8�ݜm�2�0�N�vm"�V,���r�L��u��]�Ѿ�&�\�ox�O���Vj_�|k����$	'E[�$���@<�E� ��8���H6ϕBl==���O ���I+[�LAG���s�=��;��R�	p�f\���_�k4a����bu����M��6}~M<Zo��T *L����ex���gT|<+&�v���-��(��0n���$����W��"%�'1~I��bB�ܑ��/Jb�N/h�ܭ��˿�uzˊ�uS�!0qh�i&f�"N��=��5H��K��6a��B��=����u�I�͐!��X8N�p�ȳy���!ȋ�Ȅ �
)44�&?�c���z����+�7��.�y�c�x�� ��j�����H���5vu�t��0\��\�5�_p�,4U�l�P��t
���(Y�1��{��C�S�Ab�G��5{���͑�1�r���$�'Lں$�b��s�v�a���H{y��/7R3�k���ٸ���>R,a�M�8#un�D�Ӳ)ta�-, 9�:0�����U\ܧ�:��C%���M?�$M\?i����u�˛�{wD܇-���C����giX������v�Mޑ�GC�����2%�W��m�G��XnaGiޚI&�b��2^vE&�P�r�dn�A��":�u�gJ�f���q	���q��.~��fQ���ĲTZ�r��e.Ј�LB�e��Tv�C���7��ں0���|=��s���.�.$E��T��z��vӕ~�����q�=��A��v1E��[�g��\�&�̐6	F�_���Y�Bs4{/"|�x+5��R��*�!B�4�Q��l1aP�s�>@<�����^S�gS˔�TH�cD,�'�ٙ��^��ۿ�r/;�?v%	�a��Ļ��t_�z�^�E�%����+��\��'�
1�JN�R�����Ј���o���yqWG�&� �ԥL��)7[�g���P9�k���'�ع]��6R��H؀:\VD��s�` �[D+�+ށxc_:.^�jAPƅ��$��*h܁,{� Us�W�u�-�V�~�!q����G�N��{�9	h���u�ϕW*��YHrH�m�PU�I2�}���^6��m�9��T/!����o��=�0���bb7C�����j�� u��lO�3\!��M� O3uu\g����d _��O�P
��40���&���9B�P ��w����㦃���R�|{�^Ts�qb�CF�B%z�_h��1R6�O������OH��3g���1]WPx�n�JLsH����Bs��[��/~��X ]�L��<� �0^��vk����[�3��(���R��E��}^VCYi����c����N��I�(���`߬'eX�FB������m�sm��*��ݟ+�Cʃ��uSG����S��q���_�L{�����ڸ�["�ڤg�=½=��~�Ed���J�/i�ArT�_�Z34Dθ��:e��8w,ͬj�AN��p�_.�Q�㊾6q�,s9����}�>�
KOW��v C��*Ѫ�Z1"p�KK����Xz|v�����A(qݒ���T����o" ,����r�;���$$R�T��4� o��IxD�u�2�Um��ԗX+���������fP(S�)�e=�:�P�sqK��K��vO\*���#�k>�(�X X�h�?=|��O���\<��ת8����М��.�D��fV=CS����e[��e�ӡ�	���j���b��y��[�MD2V�^�����yS��-�R�V�oS�jD$���R������q�s��	�ԉ���:0.��b�\�OK�9�Z��ؖ��'�F�R���N4}�RtS�d�.tiGS����~��v�Jf��=s;��!Y/o[�����=�l���n�C7�W#V���U��Rn�l�W�+e���(1���2�ٕw9��"���V�V%1��!ʯԚ�k�A:�%j�g��J3w�@����a�5��ް1�2/�1���g�ʹ�.�KLKl�drKg1�`詸TL�D5�M��᫺��&D�&�m�g���뜀(���L�4QJ:;!���|�F��6k�d���IF閂H �'R�p��;�#ƪD�����6#7Z67��l68�y�\��F��Y[�~W��l�)<�V�9c��3}IL�w��R��� b^"pfs���Ȳ(�j~7��XѠ7OkRydP��F-����g��Z�	��<�K+_��s��av��3'6��X-���c&�ٺ�o����ς���������'��y�\�@h5��Gp.>����lO-W諴~	A.TMWπ9M��Q�yU
�%������N�+S�g�	��$s=FH@~���(+P5���8��|U���?�_*�0n�����8$�����-@��$��@S�����}�e��ˠD;ٴ턄-{�����1��M��GtK �U��%����h�
I�M�u�\d'���3Z*`C�܁T�j�%�&��܇��Yf���;�9.$oE����gR<-�}���b���W �c*(�rE�zH�r7�팍�"y�`��,���%/���I��:zv���r���?$2�6c���h�w��=
���~|'�'P�9<��]�.�O�}7�|}����̄�v"���Y�LO�J��i�����b��lL��۰�NH/�MH�GW�>�{#�G�| �;V��.��BqA��Ͳ.\��B�%9�����*f4�8�8�!3�V���p�ӧ��HHrkI�2������҂�NCۛ_w��xW6�$�3$v�ǩ��֤�bq�%!1ŽWw���Sc��� ��n�G�#veDl�縋��P��2�/ӝ*���EQ���TH *Q���C��
�XL���@QI35)�q��,���,v���C�:����Ͽ��܃��`����8p�+�tsm�f��b֦j�D�&lS��'K��MU�ޅ�rUWk�5m&��4��-9즾�oι�H�Lzh߮�E���K���CPVu�z�JG��F4�a����,q�����'�צX=�d�?�OvCY������8ֳ�6��e�~�n��A�����M���>��v���啊��SHy�Z�̈���C��!�g�KT�<%����(��I1Զ�o����˸!�4D�f�):0�(�b�*��W(C��9��f[5��J1�p�Q��Ыk���JZ��]�g2ޚF=�<���ް��4���Eڈ��'��7{��w�D�O~���x�M[��0�囩`�>�+��"�c>W�2�v�c�k��3�J��Y�� D���Q��  �ާĦ}��\��m6�`Ӽ�V^� �1�D�g�ȳȦ��+<x�(���N���W�gKR,0�d�멏���r�mP����q��.C�z�hX{3Q!R�Ik�-�<��`��Ξ�>W��5ڤ�:��˥+��U:���pħGj&;$�#^���I��^+Nr'�����Bu������o"X[x�h�iu�8̒b�eBu.�^I�k���?[h����J0�o:��h�:D;@�S �k�9�Ci5U^�D�ӻ����R�qɆ����ܽ7��\[��a��E�^<�Rj�.�u7pٌYV���mL?�z���aw�{J%Y��_��;?f�����@˧�+���uF1O����|�g!:-X���2ESr~a����.s1Ze�k�ͬuC�^�&l���+�^���Z�X]�<���D`�X^��ћbw��{�$s��9 M�xAD��~��(���)�QJ����o�
�Ǹ0����>d�E�W8�7M��#��2idq18�)�k��(��x������V: �0 4tC\�
e9R'�{I2X��"��𑠗.���"
1�a%���Lt�/P8���p�w��@N���n(ԍ��5�ڞ0�z���3	�$D�����4���Q��҃��o���w3kC�Ó����6S����jJF/�A�ɞF��=\K�Gn�G�"%�W^Gb���]<�W ���lP��F�zs��bi��e8V~��Jt��y(����p��l�t��+���Ѷ�_�k�IS&O�� �uȦ�I{��2�Nj��LS��+���W�q�\G�J��I��99�6�{�C79��&|����������/Q�9ċԂ�!Z)m�/K�xe�8Q�%��%ҺĹ�!Wx�ʴ�
8��J�=���%���h(K(��2,J�Z������\K��4���_},u/VV��!	�G�ͬ�����8] ��f�e(��P76d�Z' R[PҪ�D�X�J'�KA�\w*���+�\�@�l�\�SϻZ�/�8b;���Y���?�����,��(�R*K�6\�79�m�Glv$i!�����5�bȿ�(��GKD�{�UQ>�1Gl����<�z�"k'����i����p%NP���j���dL�RG���[�(�oXֳ�����`�6�>��V�l*m����D��J7��2�ye
X6:L	��J;=-�b��E�'����}�t�/M F����2��z�8'�Y1w5+�\����F�|G�N�"ҩB��f*�o ��P?�/�,;y@����Vڡx�V�.�]�ZY�G���^�#P�F�pL�$oI�;Mq� eɚ>6�s�跞���B?D����@\	����P��V�Bօ;&
��8|�T�?.r��o�j�m���4N�&��R��νHO� �
7��*X�lN=�
<���'�z�
�^��$w��Sˋ��D]ڼ��P��?�,Gm�;�0��-� ;��(<Ѩ�aL�J[���^��᫳*"z'�9am�.<i��l�o&x�;s@��{X-�6G,h�}w���d���Y�O�(D��fd��v-��1����!'}�P�ۂ�2W���s4�C+"PB��Y_�`i_"}Tv5I�@<���=J%��b^F`�R��dQr�Ĭ�U��^�5�r��]IW�S���v�I��{�� &��8����v�*cD��00� T(��X>@a3�v4#���KU�<��/u�����i4��"�3&��Dm���[i�g�ތ��G��3��i0
��7L�)�М���y�!��\��Z]i��b�����v׎��ܶ���C}X�:�^N�&3�@��uawyƅ�M�*��(w�]2��YTP$+��cΖ������\������]���	V@9t���eĿ���I%�RD!���>҃����?���V��>T���vT�R����0t���#��aj��X-b��8C��X�<W�}�n� A>+�Ysj��m�Uz��$ҡa�a����l��vh`з�����X�K���u�W6
&���y���M1x�.
�� (iQh8����D%i�lxi�L�n��6qy�n��^o�<�a�qA%	�
`�e~�����:�BN�K�NP4�����^�>�EӾR�ajL�s�����S4q�Bs�&�~�g��^�<�K�T���s�/�r�����aQ��0��3M�Y�^�e;��F��v[�^���Ox���q�s�l�}�4W�/�>0�p�d����2�@r���vO(4�
�|%�mdm\�;���Ck&�z��K�55�w��]�5�AP��`���7 ަ��E.�)y%Z����Q�Ʉ]oH�h%�D<3ŉU3��<O:��C�h���3�.aJw��z�s�����<٣DpLQ}���B�k٨���+W��������y�.� �q���<)�a+�y�dC�S#V�l8� �i��To9:N	l_���_�����4S� Q������1f��ex��%ۭ	��{�IXN/��1�q�"U�E�e��˚yc"�uZJ9'h��a���x3��۔�aG�L� ��ױբ�1�[Է;D���;*C��2�WUk-fM�#U��'��:H��w:�5��29���z�%�(����dSݦ��%�%z��n��� ���6�n�dufL�	�X�?gl�O��V3E?[������4/3��:<0,�l�ʞ�/�@�NP�I�-ul�L^��=dS�Z1�to"/��)����:G1��	&Yd?��bGA����8!z)
�Ue�8�%�9#��^��Qu���Q)����/~��	A!�DN�W�bk-.�[ΑX���j�&���h�E*Ќ�W��ѦG�ĵd�	���%B�D(�O�����r\�����I��%�K�RF�*�m��b��.,h�i��MJD
4�䎴V'�mp�=<b��wP�Jw����?�l1�ķ����3�?d�9kaT
	յ~P W�ɶ�ȓ d�� It������.I��3y&2"�v2�]g������M9�L��q�!=P��8bK��O.�����d�C^�o�60� ']�P��W�WI3ީҐ�mg ^��J��[�r�3ڽ��kd(��o|�$��}%F[�1��:'��^�$S:���}��@�^Y���������&�x桅��r�T��	mDI�J������nhiw��	���9ίJe�x��ퟺ��p^F6l�b��beS '�щ������?Y,�M�4���j��
00�v5�p1�����R�։�������ҥ���@�s�Tzi6�g��b��+���ήf��;��$-,�c*�޻,�]��v��%����B�h;�c��lp��ݗ t�z�R��k����Ab4Y��I	d_��^ﰱ���F�
�n���	�8������.!��g_I��\�Z���2� ���)Cwō�*\G�.)�ֻ��k���o�GF�D:Y��ը���Ȩ�BNm��Qye���)ۯ��U�P�%қ���u���-a�,�2J.�1�:��p�m�K萲�x��F\?|��L���j"����"��6Ľ7���皎��_��}[��t��M<ν$u�����ZnrHY�/=F�k"b{%QF�&\�y���Ɉt���+�a�^���"�@���כ���vX<�����<�����K;d�@�oY��<i�W((!��$���6��I"l�b�?��g��j1��\F�"��$~�#���O=K�5�ѽ%kV�iޟ��Y����z�ϫBE�jO|��$���X�S\OM6�^�Ĺ���?����r��4��_���RK�� OO3PB�d� �|m��~��#��#(IP���ܯq�FfB��'�l�cAf��)�_�9�2�Пi���6��YZ�@�g�������+�ӕwj�'�h�7\��;�3��Cv�+)f)��TBP	R���$ϭ2�t�MUV`�#�+	��)�T���/�ȹt.?,h�L�p�Z�A�L�'Dǝ�}c���+��j�*�w�DH�Z{R3�_�Tl��o���ʡ]Y_,�5E�~E,3�2���������n7W�Dw�/�0謾��"t,8B�S;��m�z�ys�M^)�5�E��M�4�/S��^<8a���pE�Z�֭.%�ac�;:�U�
���C�ZYH��Q�Rp�i^��H�1Z����֖.u���C�ˮ_Y�ב��f�+m<[���Ԇ��lk��u��K�$(��Ї�M�		�����Z��d�@2��W�TYt�W
FhxΘ�8�Ui��#����؎շZ���i�-�1D����sZ1ąm&46�g(�WkiWU��hA�N�}��x}��@���cD�����j~�].��vzL�5y�礪 ��Ǘ��H[ۀ�o�pFYG˶ėrn:^�lY&���Oj��?��!N�t�[��N����p��w�������K��]��D>�!��#jX�&���V!w�����\$�Tm���B�U�G��D�|q�k�C�j-J�%-m�W�#�k��~���H�_Q19�-�%Z9.0~�G�YQ��*8ME\��"����Q��b�C�I�q���+�Ͷkt:�ǿ���c	S��� �_���#�'�Y�B���Q<_�.IihƼZ:�i4O�E�-�-�okp��[A�/a���)~X���z�7����^�^{?����V`E2-�ۣ	�C�����,���ղв�#���+��� ����Mf�\��a�o�{�F9[Uir�4�Md�����A��*���\ӱ'FB�2�_�S�z��PF�&�O�������g8�L&��"T<���Ys��9�P$D���ANf���bk�Y��6�l�e�;�Qz+�Q;�4���@��0y��G�\V۠�JK����݉ɻ���Բr�&L{/R}K��b����T�ԕ��"�l���?2�N�>�(�������|�汉M0�D�\<���HF����*������C��'�y?�3�ѴQ�ho�㵁�n"J� ���W�����T��=�꙼��a�}�s��ى�e6���ӕ�$l����Nh&وF�fz����L%&k��6?�sgHg�	9˴��WE0�l����t��/=��A��i��n��y�dB��1i�(�9�����Fq�Z����zӾ���!W���w݆D�3nA�,�
�R�n��^��\k��t�1n2(�r-�����Roqy�R�gO�mk�!�N�Qn��n�ٳe�_�<�
5�T�������=P�'^��(k_�m�l�ƐU�� �
S��i\Yt���K�&�L�:v�/�B�4k��}��a������L��B�R׺�q�B���n�J��џrŠj]ؒ�k�g�r����*��ﶡڶ1��+\�@�����*�V��.A��f(E����f�BB�DA�{i	��f(	�zh�A�繾���̟9��^{����O��wt��И*�wT~���?%)ģ�<��m����o�&s�_p�:w��"���)����Uq�|��'�;����Lm;�ģg}��g�t������(��3�+�P̞����9IX�8���t�![��r���/BK���U̥B�0�!�����/�_�k���l�zVZ����=�Ŗ�NV�I퍊\Nò���H�,�;>{�(�������\�����˜S�?|9���ч���lR��lz|��TWd�'���SF��E��$�N�`��w�X�ٲ��h�ڼ������[G�o�U-���	���p����b&��	��������է��X���@YC86��o9�=rټV{�'%�Е���Gw��'V-ƃO%wU�z�c$�~��?Ir�4��>����<��&�:T� n��&�Y��~h�'m�ѡ�_����8n*7����B�ê����2w�E�J�3?���e6m��Ӈ��f�N�X��ֹ��~�a�p�:��%�<�%]�D2��gb�2���I�(�[�O�o-A�m���=������ܻ�2�2���UR��?��{�I�<b]f�43+|��2�@h	�q˽��uV�!k����2���G�+N�{i�I��s�w8	:T�Z�#���r@q4y�u+���Ƅߵ>�SWu��䌜�n����t�I�;�vX�U+�ǂv�q-�agQ�L9|O�c���_ͱ�t��Q��)����F�-1��U�ڴ<�s�$T^SO1�K���&Fu��&��6��|W�}�P2�D9{V��,�f���߇w�2�2�C*�p׳^w%���,���P sUw�.);���)j�4~�t��T@Xk���Fm��0�b�����S��q�3.�ذ�M䧅�%1���"���eݾ
�T�籇���n��_��ȚR!$h��xD�lZX�	t��7L�oӬ�:�>����U��������@�՚�x�=o����ۀA�f�ӌ��C,FZ�Le��?��["\V'��	��uS�3ȔI�RS����I�ՑO	}����ɑ���³�0����C�r�%C�Ig�-[p�˵��O��)�_����U�uݪ%��
��HT�Y96|g���Ǖl�����XR%���QhA�gL�T�$D�@T�MۍȊ���=DM6�~2���/�X�Y`ʊ��	��!w)΢�[1�u��NU��I/6_�қITY׈�8��ÚT��N�ea�u�ę/�����̀��$�sF���5�)���T6���w���#������z�z<R��#�*J��靸�ǜ�����|;�6��L�_Z�YL��@26̔կw��������S{(s�žT]��{���>�j���d��D�������/�u���p{+�)��w��jn���P�^���V�������<�M����
� ���]bskQ�4Ro����u��Y��A�aj���л�5�]∇�{�FB�+1_��pp�c�c'/,�+�o	&u��^���Yʻ@=��F0<Et��J��YYI��|c��S]K3o�:��	|��֎
���ur��X�9�D0�ԃ�K���-�/q���,-�A�z�6HA
�I ����$8K�� n�n�rleI��}��_,k��U��J"�6�х>��S�a��?�)��B=�J�zVNY��cf��5��v��3�b?��Cc#ļ0HqI��L�Y�vE�N����3���ݗR��uɁ�?j&��Q]T��,^�r���v|%�\�>�о�!z���7�*�%n�gn��|�'�J(�ɛ#2���#k�{i��$p�\�ȅ���X�@�T'����l��O霈��YڰJ)��H�bOBU|��^���d�<S�vZ�K �m�q�A��u�`����C{�s^��H���N".o���b�	���+y>2o!�٦��~C���Hl��K��:;�LU�Y�[��yg�귎�;DsPM�n��D���#/��/��ۍ��=.�����?�)3S�7�3I�����k�j�xP��W�}��i�;�#��{�]�D���+�Y$���6�GWa�z���
+�����z�Ё��߹ߊ�X���_�ˌ�����f��UT҉5;T��f?RmJi�kx��/@d�r��Z�"r�z�)�U�Q�o���M_O�޲�Gk��8�^���q�C��.`oeŗ	�R3A�%'̫��d�IU�����[���ɚ���S�A�9l1*÷�Ҋ8ف�{tf���*���n���q~�:k���

H���4�&i�4�׭�~�5��-�z���.���60�'������w�45B�
�n��C{	 ���������So8��n���e9��������O�5և�ǣ3ر��7�����[��	��K���;�*�q5	�\z�j
�3��R�8��Wh]DzM�����"���8Lc�����@U����^,C:,8���$��N��*)G�j�.�4|v� �N-?�r��5r��l���[M@�E�'{[��ɾ�U�@�G��8����E���G��8���G��YQQ�� ܛB
M�/�d��V
���=d�%?
jYw|AQ�->�R��ƏU����^�Y��g|��Σx܌Zޭ�и�؟+�t@�K������m�Z|�]�
��H)����:�\�B��������v�]\k�����iʆ���-�:.kT��YX�m��*��0g���$M����2�T+��S^�&���w@��L���K9��bV��w_�j�AthH��
��uȨ/?S�S�������Ϭo�ǃsk��(�1�-�X�:�p�4/��9�<?�R�j�AD����`yS,˘}���8:����%��>���(�#�fV��).�������nN�8-D�$܏O��H����+���E4��>"�5���0V�|�r����/ٲֹ��+���a�IE98#Ut]�f�2ܣ,�ʻ��ړ)����5����0�����`*2_�`7C�]m<e���F�µ��}�p� T�y�O�1U��:ݑp?�[�_e���{�շ��M�}m<"�NG�>��I��6\�c��� �
�]r� ��e�����iE�Ʀ�gJUiEnj��R��0?��  ��ef������jK���I��#$������p� ;��X~&@8˜�1#J�fMÀȱ�V�t��	��(g�XY#����7�g�E�9ծֲ�Ψ&�����=�u̲��SNK��Y��Eɸ���R���+��M�c�z�,}�zY�W�Cy->�l�Ya��AK��"O�̦8U���X�>�Qm�%�m�<� �x�?H�]f�3O ��d��hr� Ex�]��*��Ƃr�Q�۹+ �K1�'��&=K&6���l�O!����������]��]��s't�<\�5���q�^EXҖ�)���<⧼ �	T���~��.: �q�I����S�C�ڊ�_Ǽ��ʆ�ѓ7�ZsT�'�.�3	��	�&E�rE�o�nfPl��5�c��uVz��(kR�W�t��ɡm�qIx|�q	�������=x����5D�~ sAiU��b����Q��JC��J�[f�ZAx���|�	�+$l�dW�/f�����!.��5��ˎ�~�W�0����6[/>�]�{d�7]Q}l�ܺ�1����{��Զ�Z�ﭻZ9�yAݾ�F-0������!���:����t�oZ8����������Fi4L��~��:a���Jv/�Ip��UEҌ��;�7kگ�B��m�=mV����Z����k36��W�	oXg��i��?��%�b�
�i�bf�t�1h�C����ަ�uܳ�������ț� ?ǲzV�o\eǩ���ٛ䀠��:~~�����k�&=8B���E�ԩ�=K�SwUJ{��7
=:�������5M���I˛ym~�w���f
;̬W�l��}8$-Z����N=����?秘�Y����V���_'j��C��8����ZM5���#}��z��oa�r�W<�r3<<�����eHxp�8�>:�o����z�^F�7��E��}�2bbb[����V�����m��~��G�}�":�^��թ�杪��"HZ�4V�4��'>����n;L����:����!55�]�M����:eK�szr��;��B��a�a�m�O�@HC�]��0��b�����O��4��L�)I�[k�;����qDh��pD�Tk�_�ߴ�J�,ڊ%������rd�{��pf���z�
"��5�&o �AS�/bߘ=㖙b~���bs�`�6w�i;fi����(���߽u0+xC��
}��Q�a�R�J84+��A��.<���z1��c�ώ�>��Q�x�<|�a^#�h��6�w,���y��@#��yF,~�<�QʿL]�?a��c�;и71���"�20Z�K ł/�q��,}�W���Xh�{��?	�*(X�Zp��so��#wN���ޤk�)\�!$inl|ӝ�o�����`�ֳ@/��y�>�q�'�������݈�O|���	�4�<�X�A�u	p�"���O�x���k��1 �)#0�{��a$�z���e�U���D�,)ÿ�2z������)Q���7�"�?����f��\���>�ٞ�^�sQY�>���ӕk�]���R[M�a��WNT1��$0�U/qF��8ٰ�.��b�HA�A��_�jVv���<n,czP/µ�����(K�s�/�����V'�P�nڋ|��}<F֞�ڵ���og�P޶K�g$Yo����6,.U�w����	h�pcf�ψ��,���I�b�_�>m����ʻg�PC3O����7�{,c'c/�MbSa���ċ6��{c���Ɔ�Y+%�"�i}iR�X�z[yŻƟ���a>��)�iD���9�^w�[�8QIg�ŧ'F��Ws��Y��],�bB�cHF��b��/���|M��g�S�Svs��M:n&* �7��t˱��fS|���~LQtho�Y`Q$!����a�2YN��'�(v/"]-��]�0nW���_��b�@ب�����*��"�zNuU�մ�g`��:6�7���'U%����م~�zP�[voG�x�l�_�U��R3=��� '�ki�1%�Y����:rꋾ'��}8�	ˊ;��шE���Pس?���7��3x���I���>���y���tQ��"��K� ~�.1��4���5J���?��³����J�`$lvil���"B�ǳ�Om�-b��ʁ�ZIY���y���Vn�����i��;o;��=�z�t��u�d;6�I�-zj����M�݁�@�7�<A�^����o�E�U��baY���#_Bmj}S�R���u��Z6����7NW���z���b2k��B^M�����_�k�PP�A�Db|�19�A\�E��J�n�Ix�W4�/>C~�-	9�_�Jɔ�X�B�MѸ�=+�����t�u�������z���4�-�{p�ML���G�,'Ye����[��K��|�$�={Z��%�ny��hY����R2?K\r@�7U�����E��ƐE���
�t|q�����p���O�*z���0��z�Tt���@X��%��'rߤ;��[��5�y���^���=������l3�W���5�̓_�8�w6��/C$�yE����;k,BX��e�|��0�X<�T|�>�?�	�x��I�Q%���7j8���|�m��K��5������c��WG;VY�AIͥ��j�Lש�q��,3iM�SA�a^#��R�UJ_�4Q���7��K�b\�Oc���>L�����g���'(�H5f���W�)d�߄�w�ȵ��7�Z��B������f��0��`4�ܕ������;�([U�=��<�1����l���3]���g{�5�F�i���oթ���g<N��X��P�%���.���A��b��hвq�,���?��Ԭw�j���n5�ԑ�+�\�>?����|�u�t�J����U��G}.�N� `yZ��O�Q��~S�}�g��dF��`�4�Eg��Z��Iډ,�,�U*� ͫ<5X�A4P��>|) �|���>/����R~d�eDC��@ͬ{(�
�>�ZT�.º֞��-.��ao�m@3�����0��X�@w�7Ҭ���`���5:�y�N^"f̼�V���Xȹ���p�[���x������΋-!#wa�e}���]�>�z�iÐ�N�n��1�t��"%��~��u�wb�̫���r��5�7�Z���Q(����%CCjum�����Z�h9	��AGR�Whp��u�2�8B|γb�o<���,��7y�0�� �a 4�d')�;�u�J�����r�[���8�v�Ƙ�l&���=L�R��!#Ѡ��O���Gm�ҺN�����%L��Z�RoYo��r�\����(U��kk���Q0��=4Vv��D�U��0/�!RN>3NJY�h�2-]���i�����W��0V�<�a����7j5��&"��R��j�)��s6��=��~{9����8R�A���e�ݘ��Le�N���0�C��&D4۟:���e�D�ay��Dk)(�X�gj*�Vz�ů�f�t(/~#8j��C�'�E	)��2�M+�ҭ��x��z������֣;�����*�H�V�J���4�~ 渘����w��9����R��h���Z�F��&,cdc;
��Pl��2��\H=�#��i�A�`~/ ��s�|����Se=w������v����[�J�.�č�}HI�tKj��Z����2I�p��ZvW�TN]�n�Ā����/�̛9m�؉D�XՔL9�<�o�0���:uN�}�U7�i���',Pl�_MM,SU��)Z����y@��\��/����"y�-���(���y�P�~́yu� �R<�ԀO@�u�a9沦#��Td>��{ݳST�8����>/�S/,�>ƫ�"���٘!�4��
��4���p��>En�bP�B,�у=��g|�*�9ۋ��&��/�B:����:m|�C2d���l��i9؍��	G���_�<���b��փ����1���i�P��%�ǥs��;�q�M��*�K�4�5�֒ͺZ�Cɻ�}�����Y=u��8{g4�)��~�e�mVf�g��Ҙ�Uf�(��}h�^R)�����M&G�$��m����=�ܨ�{��bT�O&�w���t�ޫ���!��÷3[�X9����E� 2��z4�s���.7��4?o��+o&�7*�8dF��+c?��I�}���A.u��p���������{�?8�È���疠?�7��f{<W���9�5��*b�i�WQ�������o�!K�V����`��
x����G0������vd���楶b"J��]���J26�A92½���C7����n6�d6Ms��)@ZK$C�ᕈ^��5�w"γi��ח�1x7_ '�ZOa�y�}+3�!���7v��r�	���=�$e���e}l=$�?�Y�����\�=��l���zf_��*b-�6�Q��q�Ѻ�n�9�2b���Lc����礓
W�F�c�$�9l�
u|�.��]R{��q|W"/)���}���.T	ٳ��#�T\��1x�4='��w�AG:{'RW-Z@�v +�j5����x���2��l��e��Y�; �bnrHu�Uv���i�
��<v;;;s���18�M2;�[�{|��2%/�U�C���-�
H��f�.�M�'.8WE�uQ7��o��2C9��gIm�~|kj�԰I�hg�75�Yyxŗ�c�*g�nw��}�9m���Y����83OXG��008� �푴A���~PY�C=�u�����_�#5�yp�}�I�� ��w ��O{�����r�_��!�hʯ�l�-����qoڪHp�"zt�̴�6Mr�e�D���2J�I�	�N����j?*���� (����a��?/�d�$�3g�02�Z��b��?��mJq�}����^����#��c2��P�h�u�qq����oE��a���W"j���ǑI��-U��K�[��O��	�ond�O�&29F	�w'ܴ
�%#�+�^���ӜIi��Ȟg�~�f	��M�T�~뗩��{ g�I>�@-�B�X�߀���o�ا�븿�n?�0L`����yϠ!���q�,P될q���3Q �����F�p߈қdK��.xNA���U�aY�Ӊ�7��w�䯫C�����i
��� u&!+�1�i�F��k�Mv �[�:�IbTT������$���ƧjV%����s��aJ��0ޢ��T��"�X�J����]�k���ˑ��b��+��=j-�,;m3���-#��[�*BS�4E�L��J�n=?��p�l�����o�����p�^d�j��
ӏ�b+kk>��'9�;�
8T	��~���2�-wT���46�p�y��4�ֆa�U�6>Rs� ��y�L���F�K��}TF�c��*��$4�_���s5m]���R��c
�>�E��: �J!�:���t�2���4�.�[��mlX�.�giߞ=-G1���6�-�U�Zco/K�+�o2H%2d���u���}����eӥ�i�%���e�H�U�<m�Ư��S��ъJ�f�ce^�?��8��t^��p��0���n$�}`ո�ʣ�T�5 Bd��:�ף���
�{7y�i'��@u��)��X�	�Z�u{�й���F�ۆ����ޡ�̿6�1X�k�KH�JH�N]�<VId~�
�
�2VϾ[�h�?��g򑼅�{yF�L��D�'d`iŀ[M�n&G�#k)�e�K������f�/��=�=�d���3��>�%X����
~f晋]�ӊҲGS����~A�H���<1�I� A����������BDB��k��%*���]Լ�[7�Q��X�i ��whi�g������g�0�C���"��]�f���2���*>ˇߌ�y��.I�T��f,�U����Oߎ�Z�W1�06�\n(e��셔R��du��1N�嶫���h���G}��X��w��q�����~�l��� {���l�5[��ہDv�Az�OnZ�f���;��W�
D���ׯ�"�2O��)~*��3�U@���|����KK��I��È��
lʫ� ��	�S��h�+�Q�X�h���$!A��&� 0��3��vY���=rN:����u+:*wY�����Q�~�I�KxE�EdݑN�ܯ���>!������#�+�q����&��oԹ�T/��1�w�����_�Ft�D^����2Y�����6�9j����%hRH	Rތh��A�/�`ۛ�ra��ZG�����=г��ExM<�y��=\����؇��%�$��w�N��d�u���ۄ{PN��b���+����Ne���
�x�{��r����}]���Ayd��?�sh�������L�\1�yL��[Sz�G��&=`���׸t,;��fɄ-�M���۩<�K�^�#Veggۉ����o��#��u��S�S�B���� 0|�W�#�ۗ���~�&�+*$��ZLj9�:4�8�!G�T�S��7ٟmB&�L
�Ǆ��8���M���RE����}]�R�lW�߮<+>"�>�yX�yd!��X���
?�c�������s�e�R��rX��Q�s��9��3w��)�E&�aQqp?���� �5#omMG4���E+���%�?D��x&0}M�d?�h6G9��
�I��%'2�j$0aHj����W�t�ϓ��0���:!|���Ԕ*Y��g>h5?�̦���Ŧ'
�:Q�εg'�"�_�,0�[�@��\>\v=�,ϑcǅ@�chB��a&X	���O�]>Թ�QK˸*V�c)Z{4�-ځ�?b�m����6���tE�BD$)�_
�hmOMi�H�1���7^�+@��Ƣ���'+yv[���$�_^�&Z���n�ݑ;/B%`�%��}��UZ��ZN��k��k�Є!k�u������Ac�9�z;EÚXD]� �}�͢����Ï����GD>��]<���-f���m(�-�)o��?��t�����C���|�34O}K23^��D�;&b�v���T��E�M�����Nf��D"�K�o�-�;k���F5C^��蠲N�2�^�8�U�H6�f�����y0K���ڰ
/թMG܁�z��&����[���d[����)����.�6Vb���AxG��YKl�W~��wH5 6��h�D�L��jV>=��( ,�z��o�MR�`i�Y�[����ad��j�HS���M2b��[�xg����Y����3)F�t����eN�ZK�%�~ �w3v�eC��?�ʞ��&�\^O؇�x�r�:X��XK��u��a���3������[ʀ �jM��K�q��F+D����|iAQn㡲�ڽw�����ɓ#�1�/Mg�O<�;Ӟ��36�c���#�߻~��_��k�s�y�ʶ7~��L��u�w�T���Tt���s��%:�Q�M=��=���Ԏ�Q�H�9��� �'�\Ȣ���Q�p@���� �_o�H�n�/"b����v��*�5��>�f��S�k�V��y�:�W-�R��_�AY��qxxxZ�(�Q�Ry�������A^�����
G�[����73�3�#���7���N�5!j�z�r�󧟣�\ K�^�eo,ӼsЙ����3R�|j��j> �uW����N�`r�+s�*�Pur���#��*1�h�]��+ a;@ݝ����7�8��h�!d'�E�@\���l���On`��^>��K�42D�z��=T 3���l·">,&�Z����&b����a�#���o��J�ť�d�\J2Uq�f��jL��3-���Xz�Q��2�[��<�C�Y����Σ�*z����ۓJ11~/1�ꌛ�r�Z� Ֆhf��*4e�h�P��Ɓu�/��C�f�B�?��o���Z|� �m��M�^��)�7ɗWuum��~9���˻��֡��vl�<l[��$�S�e�+ü4�z�ś2颕�^l�.� �U�
*C��g�9:��jh��yB_��;(����7�CP��M(s*��;� �5���L`}ZќM��|��[��4�
�����* ����_�i���/�ͯ�ٺ�a��o�~[g�(�dP��Ö��m���6�0���xc��_e�Z���|��ј��C��X�4�FJƄ�:I���S[�\�z�˝�_�����}UqAՇTtF�V�l�AF�;(V���4�uǒWP�b&�&ɡ��c�V�4����{�� m3H�VW��*�ÂR�z���VX��� ��k��׊&=�"�|4r��ׇӏ:���3�$,�N�@���#e�����W��y�s������Ҝ���q�0��<%epz���+�߈]D�\�OqU�X��3��a�QE>�+���ER}�J��9���R��B��G����c0���b|�GqV�z��]�X.�0��8��Z���U�1�o��+�˃�i��ʷ��@�����Y�㖐�o,ٰ�_"����<ǣ���*�M���,��i��	EqQ�H@WH����{X��ƓO����P�U�uum֡�ݝw� *+I��9Ľ/��A���I���i��s�v�G����Ɇ���_y���.�x�9t��\�#BV�|I��R2�������!/�7�j��G����ΠoL���������8�:�%�4 ���LH�۴��SDM,���+5ni�-��8����/(A��5����,f�3ʤ�ʪ�v�����p-��喱Yl�?��X�C�;sV���N������l�] \���&أ {(��s��j�Z�ϴYzݠ���CV�D`.�Ğ��'��8��}������$�c+�F���~�����~סwU�F�w�iC��\>Eq Qד�9+��}Yh%3�/�U��^Y�Pr'�������c��:�;*�\�0n��@�d�'�t���++b}]�?J���[���j��(YԄ���k[�w���E���%H����I~��/�������ͺ숙~�d�﨏��L�d�%6%��/�*d1'u.9�|�aFS�����)��YA����d�? ���>W�)E����t��x�~?ow���#ɳ�VÊa�`��B�������>��6�9$I;������?�뮭�����Le%wq`J�~�d�E�v�-��JN>0>�Y�W�r�[��X�~O����"����l�5#G�83k�{
�Ӣܛf�%L�?q�|����~���)<T�N�J��PG��Ki3�����!�/� �[���D3ؖ#�}HL�3�᛽X�����Q[�n_|��O��!�>�v�9�ilSb�����@��y�-fI�33l�wG�;�j�����s�?6��;�bV1��#���y(ՇRfU+LJ'^"�B��vk������B�	�$x1�uy(j�`����nce�m���a�Cf��l�ڿ���2vӠ��Zm7Z��H_qZ�P���د���3$�v.���.�SU����;�ĐrD$}cٷ&P���y*x�Lw!��rlHL��a�8��>�tM;V��͍��D��W�c'ݙ�<)�>N�jk*���%G�8�4��wR��w	l!���`dR�AW��$ʿ-&��f����2B�������o��.�����_uG���o`YC�M5=��$�z�H�.bS�sC��e��/�Ї�Q��+��+�wD����l�k����'0��C���\!��P�)v�{Һ��u�S���,�>F���}�B�� 륧k�$B +�-E������>�j�A����>Þ��a[~�����ǅ�����]s��~�5�3�UpY�xw�6�	M]o>rh�kV���:w����pu�l���Hxe"oؗe1%��P'U~��4� �
��g*�&���c��3�b%`O3��'��y~��TOl5{3���wm�s񀟯$d��*���6��*��Dx@UW�*�P}�5<�)[��1����Ow��u�]�LH8ӝ��!j�%�_��ܗ�2�`՝���tԀiv]�C6%d�K�Շ�H��zt�w���Q����7�e^�.^[\d�пEZ5�<j�����IV)�ʊ�����$�<D�-��_lB��/3{��"�0��bp"ry2+��A'���K\� �jNy��:�H+:��蔳EQ�[���T��q�n1s��rx3�\��W���o���R3`��^�~r�O��5�j�H���Wj��w_����?t{0Jh�A��+Xh��L��`1}j	��5z���'�A���#�c�d*� 'A�\�f���#b���JKP���Z��9�վ���'Z�^�/.�98�r^md������2�x�.�n�φ�������YG�G�������'�)@9�����/�@)洆�D�)*�CB<��O�d��H���	�5��ʀR'|��uZ�%^q�W��N�X��n�ⅨXt/Cg�bݢVp�[Y^t�+m�A U����1MF��&O�3��-R��Ӽt7����d�4��aZ]���U�Ȧ�B�c���{�Veo�a�H��J\ȣ����oRk��s%e�[qi�%|'�;+�3_rX�
"vGNW���|��7&%���ߤ��k=11����m��:#�������?ox�+8�/}�c�}ߒ�튉����\�*��A힇چ�s�033HW�?�%F�UZ�k��R2�t����CC�({e������e	 �}�s�Gwj�S�f<�ƭ�$~��O��]��J���B�"�ɷW�O�ϮAM��i"�sv���"�yS,��=r��s,�L{�5,*� �p�  �L^8�ԓ���,B����*_�7�4��/�3����42M|���8�8'�+9�6�%�λ�/�z�k`�7���]��J;|�S�5���A�m���������u��iR��,P�&��zR*�%"���B�kfjI[����c�'����B���<A�T�°��${ǩ#s��ܞG���3�U����1w�L�x�\��B5"�mV/G�]^�z�2����o��|�g�����si����?��z^{�B�%z��]5�+��/�iXZ�T4H&�ht���ڣ |�Y��x���,���0PG;���0r��i��2�^��l��x�Jv+�O��N)����T���<��FP`��%�o�!��&���Am��ky�%�߻l+�8H�l�
�/��Uz@c,�ư5!�8���52ɣ�����UEX��ӷ9�˭�,��M p~�4i+tకU�-]#�l)�GYQG7���Uo�>}Q 5��M9�B<�J�0�d�w�8��Ȩp4�:`x�:��j#���^�A�5��Zxe�IďjM��s�ƹ�=����x�1C���"j��dk�oӆ�j��S�������^����l?��-5B�yW����KG�5)R��r�`��XxAԜ���	�����wrN? ��YI2�����L3[�r6��V�u�?^��A�a-���R)i{2pS���f���~D�~%���
��(?V�s���wS+�����_vU���c���T.)W�q��`
)��oը���ϯA��s|�Dt
AU����%@E�J�,���U�^��39�t�HT����v��<��<؝>TD��-輄�m}��Lu=+�]�l��T�
�ɡL$�u)#EZ֎*&a ��� ���?��&�'��X���D���g�j�%��o��	_%J����D667� �� �];�=��ڜ
����/���E��VÞ�y��i���~��	�u��MлFz����W�4O�.O���eӬJ���9��b{�/hxfh��)����wp =s��c��Q���n�v�a'��)!L!����ϗ�,���Pwi��6_�dD�)�5 ?����p�X��b�R��|���!q3`o�ޅ����� ��]P������ya�X�p ������SI����u)|�c_�(�7�#������O���
��zz��(���P5(�X1�.�bU$¡'T�-�;�FE2ь�NM�$���>�UV�w"��[<s}���d�=��rW����޽�Ks��V��D��{ܕ{7�h" �ń���{%���^�r�i��>���0�Hr�JM�(�[4�\<��'�-=���=�&��h��l��aLs"���?�k��~1 z����m�*l�a1���?�醙=���n�N[�k�Y�e�"�x�U2~���O������A,��G���x;��nU�����Z��˝�峒��)�e%�l1Zܛ�Ȁ���i~7I�T�2�z7"�-� ���C�
��_蕼_�����0hU��jv�� �������g�t�Ǥ#P��󿷋(dǌ�\��rU_�P�J:�qD����'�<��H�U���%�]�TUN�`='�T� �=��0�
�K���c��6e��Q��'�N�+�J�!�c~����/�1�rd،p^���"��&�i��pcƐ�ꧡ���K􈾟=��{�@�`�Z���N��,x��������p��%������̻wr��ܹZQ����� �f��aU�K��jcL3@�̟, �U0��L�k���>�YĆgTH�w����*K�p�n�=�4$E��P�㷺l[UxFtlp 8WA���Y��-��g<e��yNd����$k��Y�ӈ𻆉�(��͡|�����v���"��ѽf������
���'ݖ[�'�I/�oз��wV�s�0��u�k�ul=Z�r�u̒���	�K�O������{�z������m޻�,���j^/���3�<�}�Y�OC�ugm�A*D3�8����q�c*kz�Я��V��r���lR�{�k���/�sa�+6�t��8ӎ���ƔR=o���o�)�0W'��q�!��<�ז�-�8�,�����;�|��P�l�g��K�❱�1]h�4ԻP�yK����>�[��/3�������Mw��I�l�D�>s������mp�޳�59������r]5uuKGG�TU���|>T�U2��ꢟ>�Ud�2Φ�����Z��l�
=�K��T�4�Э�p���x8T�w�b�&���D�\��4#B]8�Ӧ%��y�A�s5.i�n&�>mU'���5��j���'ٓ>[���j��C�{\�d���a�����#��N^AW�nvv�:��Ƥ�ώp�Ʉ�s�V\�櫛�\ѹ�w�[���_s;���Ͷ�����!��N��W�P��eb H��R�K�dd�.�T�ȕ6�Ȗjk���ՙr]z���;u��r�	�&`6��s���ɔ+Gz9?�oc���L�h6��5�W�iu���1�t�Q�:2��'��:s��>��a���r+��9�OBU�n�t��m�,����9[^.�5X��e"I���)5�;��[s=b�g�\�M��L`'��ʚ�bᜂ�~�c'-��Q#M���Cb��el���?G-y�a�E��������'^����QQv�ޤtJ���t# ) � !�"%� Ҩt
HH#��J#��H3C����u�\�,������>g����~�����w��qț����Q;����kO����[�$oo�������K���"�|K�= �$}�52%�nw���;����eec���UϜ�0�;���0�7۵�����A�����,��MT��~��"MJ�Ŵ�ʮ���S7Ѯ��9�˲)Ͽ�l"���#�:����aò�sM��fb�����ô����Pl>~��S8���63H���	������6/�:��S{v�EJZ�.o,Yf��i�#`'��|�QG$J�J�'Xc��\��d5��#���) ��K����Ff>��}� �Jz�7�X3�Gk9[�"_س�E>f��Ń����]f��𴴴\dZ�Vs܏���n>~l��,��a� ���ii���%��@��̖Z���xD�R����*"f�r�b}�-R�8��}��Q�(s�!9�)�۽��ז�8
�Ƣ��.�E��A�������>�2-H`-G�tF��($���w�|Q�tGw��+a�S޳�P˭NP������hL���Ԣ�� ��Ym�Qm4�	&))��������e�qV������#���^���с�Ч �gnVu7��ƫv�O:T)c�Q�n@,��\�fJ�H=<<$A�ÙOC�i���J���g�F���fJ�ah����u&~��x%&_���}d������s�ǣ��e���n�<Z�C�]�<��c�rE��褁��V̧�Q���pU�i��3ㅯ�$��4t�G��� /��uyN��eL�f���6"�OMuup�f�c�K��(d��<OcZ�Dٿt�44;�ҠW�/)�̄3o��T����T�^W��2q���Z�tKv��6�՗s��f}b�@i~pr�����rfaNk�]�f ��2j7ˢ�C|n�+�J%�/�4�e"�+4��-�%Pn�ʆ��7���^;T�jO�trf!_7��q��I�s`�m���ULrQ���|j�Z?F�+�0�-����+��u���[�'�9���?g�m`X�O~���z�9�w����܁9]�����s�*Sh��U���|�s�D6�)1��b�[+��>Z��b7��k5����X�9��o��k�eh���0��Pk�?��D&ઑ�$��ۡ�!�S�mmquuO<�lV��D"�ūm��UU�Oͧ� |Y�#��o�t]�F�ܛ����L���_ m����o��j1F<���+yLo��Jj�'h�_��ԧ����3z��7H�$�F?�]����^<�D=+s��'l��w��(¶S ��"��5��ȡOG$���x�@ȯ`�����>�%_��)O��c��4k�D���I�(U>�
잕�;���X��,�N˿�Z�)&��cҍY?�.P�g+���Cͻ���d����_SO/|��n�c?�tuu��^����>h6���Ԅ��ޡ��u>�WCS3��sn�=�A�Y�Q�^�-^�3vK�����@�Ufʂil�3;�����9�^V�:�N��B�}8��YT>i'��怲��A�!E�x�-&F2�f02�e�/x�
<�7��c�#���u�1�����;���>�Pbt=� �� zSXD�
�1�/��X����67�.\������nF��(��<��HWF��]��ߠ{�3a��@� 􀞞��x�bjj���9�/�y��@�nY�g�St�C�`�@jNN_��4:gL��莎�]W�*L�ြħ_>�)��`~�jÇx�9�����_S��wV�J��d�AZ7��ٞ�*���~���9��b��Kk<���q��M;��(�b��%4Z+�mt��ay�ƶ�gE�������5�N<#r*@�T��.�\1*hZ�L��UiZ>�DYZ.E�l� nĽ��M[�oib�e�ep�,�%�7��[�����M���d|q��_  <<L�-�Z��@7&��� +,Je��g367ﻸ��%�>n����Y�' iMZ|(6GrPp��GF�M"����t��]��h�g����HI���h���:Z#hF����A�G,hAY��/ "�(����f���lŵ�g����׋1�x�,��p^�%�E" ޘ{h_V�;П~k��SnI�F�O��A桄 q�v�n�+8�nL���|�飈�>��w�]u虁�3������66��L�y˞݀&605���q�����z=�1l�A>B��T��1]a�Un��z��O��F�-���#�S6Dx�����W*OВ�2YŃuٖ!b3V5*;�H�}��X?��4�����~�F�ֺ�8d�����}�S��c�ZksZ���<'ǳ.j�l'��˝�J�S���������>�r{��c������^*��r�g��ֺO�6���}"]A���3O���D�f�̓�`�吻^+}�;Nd#:Q!~�h^mF�o{J�k`h�17��I�#]c�/}�X�G)����)��?��]Ox*���x�+�C)��{{{��2�T�"�U�b�S��`�Xꅗ��\̧�;MJ�j�=�o�}>��J�1�_��{�>��*�<pd�,�e���a叝��|��$~U˿���� 	~�����b������`��қpo��^�B��%T��`�=�!"��Oaܟ%��9���Qr�|ի���ᡈ��>�7��m %hii���-'-����X��ֲ$i��o�f�rC�u�K���Zo,}�����|c��t���� ��F��CEQ�FɽI���ū����l��?�y�Z;-CstAA��ј��7Y�Zw�Ozo@��ˣ��C�J�ls~N�ƚ55�2��~��C�rys����;z���@�O�(�ڐ�� r���đ�;�E�9��Z��&i�o��Cȿ������#\gD��a���������r���wAe�k?sO�M���F���1A�t����,�JMH���Nhe���/%��Á�����ttt��<�4n'V�����Gypx8o�é�M��+�N\�z�<6C�J{,����N�A�rV�
�ɓ7y7�Ƙ8	>��*��x/SD����Ҩ�9����$Zܺ���AOi�$����=`�Vf̀Q&E��:7%H^#s���� (X���M�8Qա�;�ڢ����v;��/N����^�&f  �tG����4r�t�����f`b�`j��'���P<����s��t��7s�Е��K�r�I��vO��oZF�LUܲ�c����l$^��_nk�9l�nT,py�:�ȥ{ѝ0����\+ڨ�
p�n�~|i ��hG�e��Q��y�=��WeQ�L���g���۳?~J��}�nnL)��w]�����%�������K��P�w~/�Q�E�cZ�R5��+����^6�{�ō���~h�������$Wpct����Oԛ�����f �	O�1ȀO���� ����INIA� �D7����(n�ۘ�r`�%������H�p��Wfw����i3�+i[�7V8K���F��_�џr����h=�v���	t�l	8�ep�K��COXxE�O�G��m�;a=�@2��F���uV% �~�[��%ߗ>���c=�`VL�2���)���:��R@�A���%�γI��P�/�^>MA�#����m�*����p�V/�}ח(�?�9ܢ�����H��@�q�L)/B��cJ��0t至�}��S���w�s��v�PN��p�q�*X���=t�2�8K��l�Y��H��|���^�^D=�gߓ�����[w�ۥ:��";e���Z�k��j���K��5�z�T�f���N2~gBcsJj]�Oh� T)M�����_pnb\���-ݭ��L��y9�_̅DD��RgȖ��(U�I��9��?�)#7�aNh�$���Q'j)p����Kv{7���R4�E0�[h��<?����:�Y	�u=���voڃ�`�E��������^��MlΣ�~�]��}BV����"��~#�I��%�U��6E�#�s;�q52ɳ���yG��`E�N�����I3.��Rh��8����ӿ��j�u�B���G�<[˷,�z�<���b�;ńz�6����ɴ��2f�徴�ѐ����L�&	���M�s�g(�����bk4��ň�����m����h9aǉ`T��bum^�*���XX�2jE��C�,j�S}8x�z��NAꣃ��W+�?:ۦCͱcIb[M[D[�����&5��j^����|�Y����7���	����򙥚�������b����b+���?���i�d�>��������>\����*��4����1��/ƃ��]s����\�1�����O� 	neoO@DDtv
sAF�_a���S���ښ߲�����Kk ���םD���_O�]��kQcHB�������o��\�>�]�uchb�6v9�r�=���`gh;lv!�Ȟ�i���������.�M�,!M��j$�"��;��l��j��^m�r�v��W�/뙮�����S<i�@���O:9�ϾȪ���Y��6?�9Io��u<ʬ4;���<��I����� �c'��ߗ%���o�<�n�71�ۥ53%���A��pX���ry��xԫ�]���4	{,]W���'�ª6�L��ʼ�
�^�����5���0�@]�87���Ah�ǁHP��5���M:���y�(�v�m(_�.��I-���gE��6�2���w����MЋ��vpg�>4)}����i�MK�S��fg�ox�+��kvN���>�D�ܙ���E��:�����3�U����w|p�S�l�8�7,��\��)�uF�?)DHOQ��N��((���oֱ !��	� ��l�To*���$�ഽ��v��7��-���=Q��Z1�����P��}ޞ���$�Dm�ry���8n�\�Ϣ?��%���{�������Sy��"��*��Ȍ9l�%>=�t�<c ���\ox��:�������S�r+ƪ�>,�zB���g�.G�ss}yvs��4����O�a�ێ6l������4�z�T��>48��oӢ/�옂�`�~��<yA���`�mgC5�;! %!	h����X�G���}�� &G������������e.6lm(-��dI�������^�0��c����uO����tbYe%��.�ٿY�u�N JK���f{d&��!ٹ?A�Tvd{X�_f�M�������/��6��cjhW�||#�)#���`o��-����V3"�55��)���hU�Ԩ�fF�cnݐ�MG�Ю����V�ǩ���?>�=�yJ���5Ɔ.dd@P'Mz�#/3�s�;�������W���=��3��%	b3QOڭOV|��4�^dț�i�"�q�,�������Ht�1Q�y^�M@]ԏ�����M�IK�E���=�M'<�<�	�~Zi����1�gs�L*��� B~ڍ�d���#QMMM��.����=neee��b�;�+�-��5���OK��Ùە
��W����hB�>CJ�wW��
���-�t3]�	������Q�zf���{LWm���ee��}t��}p��'9^�����@�W���N~��g(Dk�j�]�����]��W-7�,��⻊=Z<�����떖������E~�������#������c�LXO���� 0us����=�~KUU���5`7�I�T�rc����;��y��&���m��w������R ���Xy�G#�(��ió4�A���c���x�f1��Q�tKU�^䞴IVM�7� әL���1�K��ǺW�Y=����wa��G�e�I�ʪ�Q�sjm�vn��:uD����I�O1qh�p30�Y\��)C�! LЮ����x����g����	�o1���n9���Y��� ZP���g����Scs(x����"��-&��-�7�u6�����k�h���G�1�ЈH�,��!����s$_}q�}w�Ҕ*?�����^�zD��+J�������@���O���ݲ;�+}(��\�����!~��!���zB�k�Jp�S�o�L���Qd�U���Z�*���=�S��f����L@�W��4�w�_��-�`�����j��Òq�h-�Ǉ�u3,�{Ⱦ�w��r��q����޾I�AO!�M�Jr�%C�D�?���_�-��� ;<�7��%���NH��=]N�����8x���c���ؤ?fXnoq������Qߚ��gU���L5N��7��\����6A'�Qu��x���9�w��F0]��oZ���:Z�̇�U�D
�T�o�(��w[�gp�@��ΰ��9҇
���#���.�'4w�s2e����=2b�-�^S:Y'��/�Jg��7l.�cuɞ�kP
U���s��N[~�:֏�}������1�T�y$�o���_�l[��f�KZ��ze�6�[	~�Sc;R�4h���@�����L�o�R�p��/�`����eHN��;�ݐ�C<w/eCC�ik��Y.�M�6��,�!�Ŋu�J��ٶ؟���G������~H\t*�_Q���ґ��n�R>��!�h�Od�W����^�\��| 9y'N�����F�Zb��U`�i�(�b�Φ�T�������_��my���&|P`�M�P�K�*v善�yź�er��&��9���}`��z�?�!�XhqĶQ�fc ��Лr=<+��U��
����Ϲ��N-�M�+��-�y��/��}�����ѫi���5It7�(' 
г́W�uF��U�q����#�,��L[����e�%���NP�'֖�.���FKԷ�͋2E��O^���z���XI���T���GL΍�&^���yէ/,A�z����ux�eAv�$����{Ƨ���"�~=)ƱE$�/�� ��|�(2&oo�������y~o$[V�%��2�%��A����[DOI�@��8����j�H� !��C�a$Kn-r��-�t`�.Y+�_��� ��������ȘC�;Nv%@!�o(ۯ�11DEE}.��ai���R7oeV���њ��Y�ou���ߵ�v�����Ԇ����o��-����k�5�Z�F��#�����g�[P��{ň5�u��� �v#Ka��L%������њ������r�痊v�	B�.6h
�WK�Q�`�9�-����8�D	6�|���@���_mH�w��Q��2����ƈ����ux��e�E1���K6 A7+7�skq�f�����)o�._^�1ږb�l�4����AK�z�`���0�rn1Q���r��)J=Օ��l=KM��&m��!��b������	$�.I���QXT�1���w�i���V�j��x��B��rR*�'z.��H�9��U@�`lQՐ!8wKWՔ�$cN�+��'�uƨa��ɝ����m�ݚگ�.H@Į}Ք똚�Cgv��C�㱗g[����f���^�1_S�^{]���dw��5W��_��)���#������[��xv��T�-&7VT�Qlz4�]f�vA�J��{Ԯ�G݀];��<q�u3@����!���U����:Me}����C�B�l�����J�!ᛂl����G!*�(�fe#*��{~��U�(�����Ct����� �HH�k��"a�B33�������0��m���ɼ��Cd�gJ:<�kP[n�����.�!e�y���3�!� �}tg�8F����%*��b�����7�zfO�]�cM�>�-���ϩ:-8a���~���CԦn�1�f�*��z������p'?�ۀ�Ҡ���oNѷ2 >�)�zoQ�;�ēT2"J����|���\^b`��Yf��J����7�5:r������*+��+�F�R�t�_a߬0�`��&��|�!1�3���!�,��n����G�o���V���\�{\`hi�k�q�K�!Ѫ����j��:"j3�BT����cv^�.8�H�ǌ������,���$j���[[���������|<r����Cd��ZE�u뽚�`��/���}'�)�a>��s��v�����O���ؖ���U��ꎠ��z����N����b��_���J��"�J�W����m�)�X~��z��a1,��[|Z��-Z~�P�̿9Y��ߪ�Ř���P]�R��������X�3iV���{3���āWk������o�))uW�X��ࠗDd$:꼠��O̬�u=<U׉u�d��Meϛ�&�H��T�2Ƞ� _�ۉ8�MU��*���#�����M�E>��Zܶ����I�5���G����E"�3��c�]��iJ2�o���2?ӟ�\E��ߦ�q1O�x?Auv=�q�U�dUעd�G��\�r��/����M���5i^9^�ݟ��Q�̖ `mq{s��E�o<d��3ݑ����f~H�� �I�����*�sw���9��$�O�x?Ӛ�;�S���pU0�J�q��j����O@rm�$�J�8/m8�����Q�i�|G;#�L���r�� F&����Tw�Ӝ[|����}��lH��
6'k�\�p9ܷ��U� ��O'��c$N��'��Qc=5�(txS%�A�X�E-��`.}Ukn��-���ڪ�)r�~u��C����ׁ�����ؿ�b��x���>-�����KA�����q��.�+�����)��U1��Sm�q)��;�����4;�\��d�a%�Z�O�hꊒ�֗�Lx8(*�qkQ�R�2aΙ�>n��I��ק���*�r��S�����+Vt�b��� ,0�R�s��b��ѱ;3i���+�'�]B���� �F����?�M�W�E!�~������֜�8���,8+=X�P���L����&=M�j�^�
c��I��d�t�[C<w�H��g�僕��[�z�����x����ߋ�����HI���^�v�7To��#\%������SD>�1�5�hee���*w�Cs������?����d:�ު�W%6M��g~��ڢ޹��9�<�8������W�j^\��)8���G+X�����H"��ܶy��B-��rEz�WL�	�,/6��9�R�rM�_��� X�/�^�:n�j����	��7.j:W��w��`~��f��'��[-��������?���������(+4e�8mgV�~GCm~O+�.T�w���a~�%O���G���ˬ�Rߪ�N����3��̇��z����dy��&�k����I��FF��IŜ�)S����)����.ϵQ0����`��f�ă�����?m�}�S�uj"i݋�����؟`"�'D�5�1�$��<:�^�( E����t�d�����b��b�5f��Mt�������t(�P�=X��)���	6�����T�=S�����إ&�
),|lx}�xs�[m�C8����3���C
�Vf��jU�M��[���`�sm��r��b7�*�>�_�EY^���w�7�nj|�Nl{X���N��i!�ǟ�����s��@Q��F�[�f�`�e��b'��L�P',�LS�R#��)�"�����]{V!d� !���_-��+:cF���u���e:��Ԝ�ِB��s��@���'�f�^��J��ճ8?\G��/�/ ޛ���I)�OX������N�����^x�-��G��(��O��@�X�����ß���f-r�o�`�'��<�+����8���W��Y0���u0WT��%��ή8�f�4>WR�������ä,Kه3�ey��F?&��(�JwB�I<g�Ti#_=��Rt�Tx��v$�'�Q��	&��������P]h�����P=��~���?N��I}�X��5̻���J�f�V,r�l�1B��yx,	-$ ��'d��N�$�y�/n���3l�	�M_�M���,�ݼ�B1�W��'����D�.���p���T�C���>���J!�C�v���S��(�Ɍ��7��w�2��u�5&��Z�!?T	���;Bg� A ����[�(?i��Ӣ)����Z����s�:�	h��0�c��~��&���zc�<ztn�C<zi�����c��h*��3�'���/:x���T؅D'�F��Oʹ���E��^E�,N��*=�F��p��k���^�.2�݁�V³(��oS�ܶ���A1!wi����1�=c��x�j�:�C�Z��x�^��������9a=x����A���X��^7���#g
����0=�	�H^Ϲ���ִ�SN�M"�����G3*�Ot�L���E���!�x��������S�z*�A�bl@��a�-gb(Ѭ8�Lp��ޠi#=��B����_Qe�3���#��,.�`TŃCD:�!�|��(��o3K�W�>\}+���K�G��+���_���B�tO�Y[���������B�Z.�p��o�yƂ�M�����WxC��"���xB�49��W�W��<	mEn�����c9=<�u
bQ�����s󌸼�v��n�%�*���E@�����̋�D���co[
pCX,��=�����=#k@'zeWT�!p�� ��܎3//�y1.��&��Yl��m�Q���oi����ʳ���߰�UN�#����bhi>���_�V�f_���Y�U�t]� e�2�9Li��9P@`�A5V�Y7��Q�����O��W��Ab >)�h{�8|^�g����Q6ч��n��f�lY�Y��IIP����d(�fe��P����W1��3/��y��o��rx���apOQF�{�D�ë̇���Do�����N62\���I����g�kS��ëv^�*3n /T[�1��%�D<IUQ�D<�9��!م�Te{�%�CĽ	`�o����hR(}�B�����&�
���0q`b�×�"��ԃ.����#
�?��/�ݨ4.��"o�B�4���^���2�:�Y�1�|խ�6�B�/�lE�˸�┲|�~D���{�Q� �(����lO�ݙZ���Ns�I���یc����*�~N"�z�=�sj\O6�"���=��l�9����T������s�w�o`aV������ �R9cD�a]��)�n��y�L"d�����&_:�8���h�N@{���Yp�f��ч�l��(�Z6��'��3�:�N���(�Zh�K���A�t�j	 �)edḽJ�X�(���16?�&j�
�n����Ҋf�<.������N]~�\�u�##�`q��61J�܈.��I:|VY�-t�!��c&R/$Ȁ�y���:�'-�<������B�XxF��$^���_,]]�?)�W�w� �e|�l�xӃ���}��	�I��Um4�U�LC����߄�H
��S��D�;�u	ݫ����@:g��[KII���� ������`	���ѭ�����_��U1F��J�0@��)狰��|�E�:e	��Df��v�����������E���]�&�e�mMCj����d]�"�.=�mᘘ ����N-1�YHԛ������vG��w��|�SE]os97���z}m����sP(��f����yU��䫲���>7�H��Y,��6K�6����V�����u\Fi韏��4h2F���C_y��gzD�k��K(R6j9@2�/�����}�A���͵�%����g��XIrb$i��{���u�;9�b�����{%�%\�"���1Z�M�ۊ���� 	��� b�XQ\�Q�/��͐�[��j�H��U_<�e*�����+++�\گ��]c��A��!:�������쏄���O����-�E�bh�.4�8�W�>��m��=���'�����c��L]}�|�_�"�<o�/�8��J5���&",�H����:�E��@A�'tP�	Ff�}����+��J O���p�[���4/q���	]7�3aq9��"T�g%��d�9�_���q��R@�چ���^t��ϸ��z���K��i"��l��q���%�8B�yYZ�C0��������B�{���Q�O����bp�(�p=�u ?�Xd b!fIf0=H"׾�aW� ����љ�=v]�PW���ʤ��� ����$}�;,��<�ʕ.���*'	�XL	�T�*���|�T2f�T;�����ڂ:f��Av�N#��s��_@[�M�m��<���*8Pox'�U�4}����O^=���Y�{��}́)�}��Q0�vƓ��4�Io9K������<�"Zm�#kV@
�?y���矼�AT<J}˭wjH5�ҙ�-����ᒬ�8��ae�ǣ�B]�ʓ��R��K��Uy|�����"D6�fsW���g��j����%�?C4V��P�&��ԥ�Q:�O}�@G��}%�K�m��b~x3�nl7���MqG��i��H"H;s�"Jͯ	я��F?�O>l.��<^~28�]���"K��y<2�t�к?\t���Gz��mY�ٚ��R����/+�s� ���n���!1�!�̋�}�5��D��}�o�4Xib�f����)��B��*�� b�$�
2<�3�_�Nt�d5u�e�����3���="��sOW-w�%ۅ�g�s�(�mn�tSw���������x�i�J99iD�����-t�~s�95��I��:\pRs��XK:�w�T��2��6lyJ�vt��K/�
���+�/�����/�|Nb�o|�'wO?d���"�C�=W_Ա�jpt�r��[7��Di�����eaP	ٴ�T�V���2�jD�??�i�LU��Ej����?�����t���Q}�We����%��@ �xcw8	����X�\dJ(J�cs�����h~,-�r���r\�~ɍB�'FK`�gK�A������T�h��`��-'X��(���\�
�n!�)��餪�V�QV0x׭����R(}u+��������o�wR�_TD$���FIw-�0����-�«��W�9p�Y����ӉZ�c� hP�����5ml��T�ת��v��p,��z��l��&djJ���]Ĥ�yMMtCCC��'�o9Ҹ#-Y�8�����3��)�k%�lm�B��n���))5� v~�Wݖ;�0Z��OʉE9}^a��䎚*|�Ӟ���z\Cq�N?�X���Ċ��y�+�Ԓ�hP1)���o}�b���h�m�<�z�Ѽ�F"���O��|�q���&:�m��#��o������]*�ݒdz�O>P��魂Vg�μ�w}�~\j��d���:v�s͕ţ��H�A�*c��?Y	HՁo1�sBx�^���c����M�x�������:�"BBA�x�,L�׭���Y�'�����r5�B�Q����8w�_}�r���́_u���z�mN̥�{D�ſȟi��$=e���I@v!��ܮ��dN&ޢ՜�fȪ'����m�\�
�Tl���nu�?�tY%p�g4��0}~����� �R��[*ܦ�\&w��7a�����e�GO�f�c�48��+�>��?0�Ls�*aـ��u�,��+ޛ6�Y�4���d��7p%���¨~�������	�zKr0M�ރ��]K��CRF)�R�
����?��4�O�o�9������o�n��n ��!�9D�+4��4�)��G#�a:�I���	�r�H"��S|=�@z=��h}cv.R�؇r�0�1��I�k������0��M��*�������������)�M��J�er#����bI�&���#�ϋS����K�b+�{Q#_ԫ��\w9|����w�0�V�d�wުW��@�j]0��7������&��oV�xk�4�u����_�I%h�_"Y��0w���~�m��b!�K��1C��+��e`�3���E����|�	��5��EP�B�ʷ�b�`v�������H"�H2�p�p!>�S���~��z[��X�©ߊ7حd�W]Be���u�7�T#�Xs��X#��
i�Vc%��a�\�X�Vթp������?���Tx־�P�?i� 9��9�'�����/�
����ޥa)�G!,ϒmF�P?���$�,]@�y�+�eQ󡽽/0����-�<�l~��g���57�q�s���={hm�}�`}Iz�q��#4"�K�������T��0��u����/ة�}~&�V��N9qs\��oq~��~D�X�.Ǯ���A�kĒ�*������&�V�;�:#�cTr4���܍���ɧp{/����e�УR�Z��h\����7k|0�ü�A�H+k�z���S��ܦjbX�S�KK�����X}\���|.�T?=M����N��o a��@�7�&''Yi�}O=6�Qf#]>�t0V|,��+�y��>�������18!?��Nӵ���d��n���ɮ����2�Gy1��۝�d�t�m��}���s0+���v�/A��}B�mx��JZV��Jr��$i�W�9�u�,��K\��$�L4���bD�Q�,}�Y���E��;��¬l���Ȓ�I����NLFc2���c~g�B��ɿuuu�0�l�{����_L��͆x;~T.��NON��lc	n�*<����\��v��{�G�[��<Wko�����w�`������Eد<l.:��GjO��J����o5q!�m��;~V�;��/�ޤM��G8��#qv�3�<,KE�ȰC&����?Yu|?D�'#R�����Wq#�c!�� ��f��T�a0�W�0�$�)vf9�:ڕQ��6�� p�+���@�&7�5?O���H#Z��WGe��|���؅�lC�n^__ch3��1b�/�.!PEO�\�l�ͷ5��E+o��tf·�"6��P��|��5���3��}�:Z�>uͱ?�|s�:���|���E���)fg�<��W_�z�L���	��'�,�	Z�sף��.�`߻�#"ʈ��!���0�~.m�9�ß!y�c�^m����~Չ�xO�=Q�Z銨���r:瘍�
`4�ߥ�x��1z�����H�xT�l�V��w�k���ZO!akgf�A_է.՛\��'e�B�9^8��b�l:���U����M]�Bm�p��*����^�
e)�o�ȹo&�~
Wj�g�K�h��[�z����aP��Q�@m_��"͜��I�fi��w��	z��t\ ��#q�y��)��+"�x�V|*@�;��~	>�iY%�[%����ͩ�7�NՏ�k�3��hk�;U�5�%�5dv����N�b�737'���`U�wed�m�>��e�m��rs���ZT�'�v��n����Z�%�M���u����c���u��&�z�,�:6�.a��8�nاD�JL-e�uև���/¹+����̷�r��h�غ���C�j	=�Nt��]�ga�ں�v\�Y���.�骎C�GՂ��3q-����G%lI��S�
Y�4�ۧ;�&%�Ƣ\5�I�.���<З\�ڣ� D���ZO��� FD�iN#�"_5͘_�$u���(����0���\T�G�lX�+�p�/Ow�Yņ��s\��"��|�G�/���Y�"x*����j�>|���Ŏ�@�Ȃq��I� �W�o@�������+�~w�� �i�7�%7�A������"�]ވfM��\�>�3�Ưg����ZIz�J{�Rأ��g|�4�UQ!���Vz�2n0�)WT���������P����/�ƃN"�D*I�!���DX�����m%��eX��Z��� ͻ�ܓ%s�%�u��d�u����|��!��aј5�jF���}�E��H�U��^5���i��UY������%%�L����P������'�x��8�� Ɖ��ts���1}�'T�E���Y|���͌\#��I]ގS ����g����E��-�� [u��ۈVl ��}7NN��1|�'���,�}I4L$j�J�����>mM���ʋ�����B'�T�ah����`�$���_���^o4#/�g׀#�~�A"�n�~,1�2r}"`m��fŒ:|�
Zb9�>_85�+S(���#\��0퍝`�pVT��%�w��
��)H�H�w���ZT����Z�Ԣ�]���sV��yGϠ�������"cX�%�SEf<��ۈ�M���ܟ1���|}�]�B��Ƿ��>��}HKf�@�cNW�o����E�������#�ǆe�΄�*�b���^δ�% a费��:
=ܿ Vd�����(��h��H�qY��nYW�� ���L6��P�I���9q@~bs-!xm���*�e�Ͳ���~z�����7%�ۛ���o?�6��=�o5��2�0���O�>�|�� 2�b��1u���W��w�m~����LC�?���Q)+��r��|���\�f v�$����������>��֍9�6�v2#�?�sv�-�l�ڭ����`�7���|Id3I������z�kGߗ��]��7����G���Y��K8�#ސ� �@Q��y�	S#{p�O^>�!$��r��\<�I �U�������Q� ��T��1�r�̀���f��,,*)�	D��۷yVU^������C�
�� ���������ڹ���2}�c�����V��	y�W��k�&��4���j'�x��ဤ�r�m��">�; �-t.h���c�#G����; �*���Wb��ϊ*�c��?��#��G�u,/`>-H�1O:
�(�9��(E4,~e%�h��z���X��B��l���%�#,��+�Jņ�f���8�� ��ԩVV5��
ִ�V��p���_�2�\Q�ٸ��Q�=�򱺥z+ ����f:�)p�����|�eTUa6Lw�$�i�n�C$�Cww
�ҍ�HHw�R���Cá}��y�o����u����{f�k�����e��u��y�(��<��d�X��Np�[�E��T�d	����?��{����dƮR�q��S�\`@4�|m_��ל����=��6�S�'ϰ<S
-��h�<:2-�%�>��Yu��?Q�������qw�i���q��_ՙ�S1�j�e^���%Ӻѷ�D��9M.�P����}��ul��FX�\�����GGO�V��,̟|�HS�ϡ*�Z�2tL�<��'�}���_�����5T$��E����'��[n���i_�o��9�h��<�k�6�3<��6U�%5O<¨[V��s &�<�`/\
�i�b��� `��J�߆�K��$X����y�fo��7ƿ/���n6Zs4�3�6b���Z�Y�+6�Ǵ\�C겋���umC��0Ye
�镯9t���я�tg���k���|:��]]��JA�t�LYbf��n�����W�㓓h^y_�����BqN7�*7�0ާ7V�X���V��T0{:����a���	�D����dm�wc��%�7�U��їgU�	�
��p^�~<%b��7Kx�x��_'���{��U�)�X3M./��x]��ml��W~�՞�[e'<焾��e�dB|�|�����*1 &x<%$�]	)���|ݴ�AZN���t��)����?Z 5�����묢��8��0�DfX�!���kV	��SQN���A<3��"8��5L5�-1�|�b�^Hw�,e��3�l�c �q9'RNx'�
u���X����{Eϰ�J�a�h����.�ϔc��EVJ?uCGiIJܘ2���3Ѷs�ul���M���%����\�=B~U�� ��@V��B�wM� �P|ن�����&hy??�� e,Ff�.�u�<W�ܦ/OR:bY���xqY��3|�o���5��b��d��'��M�rmP�d��>M&@-Ԑ�I�G�|w����~p�YKpӄO,|g5��TA"A��y|y�!L���k�f<�.�͗y���gz�w�����n����.K
�j�n�9�kf�7r�Q$����C�O��φ<�(�3C!f0�헺L�2��R��}ۓ�o>�0˜d��֗H,�� ,��?!PYE5$�3������js�6�ߔ0v��~<��Ҵ/��r������i�1DU��T�Ř�#�zBB�F�o��gRBn������ƽJ�Ӛ>�'9��Fq�'�ѴC�˼���ׅ*�>�!����O�+2&Î'��<�ܤ(>{���r�V��,�q��"�>��Ņ��`[�D��7!���ϓ֬�F��/)�����l?��g�}N��v�K���]eP]��GP�q�~ܶ�I���M�X�c�6�Rŏ�(����Ē�����)q'�Ii��X��ؓh	��D��W���~�F{w���W2?䙂vĻ���z�Z�������V0�!��C��*�u���J����za3��}�����N\��&'�����*|6)��<i�V�2�"�bA�&�?8�� �BW���~lm�+�\6��o2��V���1�<����/�o~繯��|�+��,����R��g���h�	L�\7����8�s�?o7���|��� �+�`��JZ����.�Cm>��/���kI>�n�߳�7�������Dp4�/�^h٠�� .Aclhjv*u�K0N(A?�5��2�u����Ӝ��J�zfJ�vhZ���f�iZ��nyC}z�����^��Pf-�w����1���m��b0j�K��������t���v��{ގe��w�	7��4Ьȼ
߆�OOs����	���n���M5�@�=?3Y�ӭ�&������kc 8<r��*�(:����Bvp��*�
7��혉�4����ަ!oX�is�Q�\�ا���n� t.��Ǟ.����z2�u�V{�Q���X�i����M��=�����,GD����d��PB�f��s'/��v�crjj��l�P{��������w�U����2��NF�1��Y)L_t?�69[ȕ;�`aDQ��:��G�^�����S��U�ݣ�*��P��dY��G>9��}�����>X/O�����͛����Tv� =�7�}o$]廃���W�B��w7��Y��> �|�n ��f�{
���v���������8aݞ������z=��0���b[�\�W}�1��b��L���_�߳k����QҐ��n����sb���X� Ot�^59����#]�T���߮�k'�|.[�uF���]u|����Ng�����Q�̕�},Ƥ��>&�������e�#�>�E�3*�^�-.|����/��6h�������OK�_���K�':�8���p�nڨ����Q�z�(�h)����!g�$+1ƷL�o�5�rot/ ��'[-�S���2Ja��y�<���XW�V���^�x��҇��q$�d� �=j4�|��-��|h=����c�����kjhl;d����CS��g"��D�_�/G�4=���j/�X0�(G^r��]5<l��~I�#�P�ipEiL�����'Q����/
2LM�����%_��C��OG�4����+��B����TM����P����_�p�a��!5�>�N�W�⿖��4@�.�󫈛j����Sm��?N�GQ._~�kyĲ�����p9Sd��N��?�U>]g��	E�(��dJ6$,��ǫ���/�m	#*Ar2����r%^����B���Ɍ>U�>)�Nr��� p�L�N�{��lrɖ*�����2 @
��d�F�qu����'{(���Y{ZW[�rL zr���b��t����:�D�"����t/л ,s`�6�#&�+=
φ��D�'ïuy){��0}��, ��WP��@��?wn9y�?�#8���/4� $M���{�/歎���eH����?�)��7x�޽�o���g�	O���z���+��S���䁐q
D݇wE�0x��NBp�!E�Y�O�c�N}:�E1�g�$��m�1͸5�
ޤ�Y���7.��Wl��&����W���D����������z�5	�c�m��1g�c}zi~>�~��t���ѕ/��{���Vo�D�K+����',z}�v?o��,bwdќ�N�Y=x4ǮI�le�4�5�~�����C��֏���11����;�s~����"��|n��J�� ed%�Sâ$/yO9n=y~ZF�X\I�齗k+�4-2!W$�´�A�V�G*~5�,cY��ݙ���{�*ġX�~�+�����G��3D\�P3�����/�$_'��#"8��q��� �i��ܰ� �1</@�VMc��~T��g��jy����'���g;Pa���Y��%�Z >30<��i5�����!kK���MUt�<�
�]������9�h��}
נW�8��qҖＫr�:�#5�Xb����pV�U?5i�ʔ,��e��c�y?�����}�ȉz�רZ�'�2ؒ��?S�
�BZ��w��q�߮�-U�(F�+aӶ�E��5&�����|��l~�M�Ǫ�vz�<ն���&��3>��
"��������D��p�a,v����iA|999p=_�/�B�,��- Ɏz����k����O\�ݧ��(����&�t�C5�A��%9fb\ae�d�������-�R���r���ѥ<:O�V�u��N�z"��}�	�*��bλQ:�.�����`ko����u> �s��u[�[�׏l��wg�MM�x��O{���YV���ވ��SfYw�P.�
�v�w�)њ-�ּ�z� �X9f"�:� Gc6��N�T��Z�-S��b_֠Aj;v��h�?�bH�B)D�`f�u�p���M���PT�D:DM1�7>(�z@��kX9�76�wjD?o������ԧkP�HxJZ�zݫ�%|w��g(S��O������x�}
4��#,|��@�`F��h�YW6"����Q:_�ji�!�ó54��l��;[�e5�j]<...��#S<<<�}�"9b�.f�]�#D�������1����(�O���OY������ƯS��7麸�u�6��#������S��)���F���Q�Ϟ��U����&�L;�̼u�/:^㼱y���jX7 ��,�X}�m�}����$�;��jm�X�s�8�����ln��'nSv^V@����vӧ��l��;Z�B+%���R��z���rX��C�����7��%���,��x�>Z�Y����A�bWۗ���2j]������k��rzw'�޸������x�\=�d˧F�3�s[t�tg�q���9n�,q����D��:�����M�l�_W�#�:��<��ӴD霹P��`2�u||iyYE�n�sI��Q2����H�+���:�nc{P��~RB0�w�<2=;?��?�U@'��s�m ��'ͦ���XQB �MTj�y���<;�s=��k���Ч��sP���v��%/���)�.ki��-��>��r��WZx��
Q0N�����=��J���zF��hԞ�|��ۭ����^@�6����O��a.��Ŭ��c1���{0;u�e�,���5����$���	��䋋�T;��n�]&-�*	�L�����ځ-�j\Ѫu�*�� @^��_�:��P�����I�xv�>Z���Ug2�l�f����/��Vu2�[8)�ql5����8XX��s?֤Bcj9կ�6s߆e��|�_��;������[�BH�Ȅ���!���e;�~��O&ޚ�;Y��c�����/?��퀯���{���Ѹ"����t@@�¿l�~ߙ�����i�P�ceXJ��$>K� �,~v�T������\�Nt5�m,�0��f���q"z,��X�K��J�y@���`��!�J����Aw���6��tt��,�j�Ƈ�ŋ�r�[i���zE�EnRw��P�D��=�����!_I�d"��T���""�<#��WBN��=Q�eN��X���YX̴7�}�@�*li��FQ�#��7Z�o���#��W�-�u,�S����D
�<�g�no��`�.�2�5���{R�T�V�~��9 �Pf��3B�L�}zz��qjq��p�>auJ�=����w8^�6�!�+8o���K��(Q��ag}R��hk���c�`Ϟ`�^�� ��Q>$0�*�>���:1AQ�W�q}}�x2�/>6��������8yT��୭���,<||��Ck2zUY�[��<U,F�q	�導��Ƴ��lܰ�.���RX��Y��<��`y*�RV���%��}"�D�׺�|��R�b���qcXl�-���k�w�bqryMMT@�;�,4�9QX��D��/��}��t�@m���˼O��s���&TP.oL)�a�C�;��h,�~�6�Fu
���&�.�/�O)�����؍��$�D_��cK�`���4S+0��y��Uf��Q���h�l���$�҅rĽ��uR�w���|B���lu�;�^.{@�p;�:E�?���i��V�ߌx�U�1������I��1�j�!�)�]�3���YP���#I�j��eNV��7�#�h��Ԏ�|���5��h�t����$�(a�u��Ky����`_SK�ʊMTL��r������p��r��lи,�_����F����YX|��87UU��Xk�gՌ����Ja�f��|���סMKy�������aT<�V�T�L�̞2ΏB�?���[���{�%�w��S`"*7��Y<��J� ��ayy����6y��/�)�ttt������:M�A/H}��G�T�����aU�x�*!C��X����
~-��pՄ�V�20d+�@O�Q\�M���C=�A��D�&�H(�&r Q�˽C�|��NH��7Yx�I�F�D��k�v��ז4���IDŭP}ʲ7x���`w7;��K��S��H"��|x#���N����$p[�o������b]�"N[Q?���Ґa�z����"���Taʜ!H.�[~�6Z��P�c�>5��m��E�Vu�5r�8����C���9o�����t�p���,���Z�>|�Lk���T+N������ؾ{SW � W�Sq��7�`[���6��r����N#n�ԱAඬ�`��.V��ÚĮ��>��g ڃ2~��f�U��lB�iM~�(<~`�#���<Ԡ��+A�C�
�2~�st���f,r�a�=gDi||m�f�;(Ң;F�f�=�~�K�9|5ۼ�Fb��Q�(������3K*�X��&���[�%˟g���U��#�-Ǜ���.w�R[�W�H座&��===��n����Z���Q���;t|��Xi�9��/�䲍�h���~���w���>%e�:8�ޤ��"a���S�
�u��5���WGK{gUXD��%��/�=z�M	i9Vҙ���P	ƻ�\A�搰n�k�>3k�rhXߤ���������;�V�*	F�����<���iI�䪢"�Uf�[OmV�1��k+%��Ye8��ȅ,������g�T�Uϝ��\�ŕ���f�:-(�s��(y�jN|������O�UΛ�b�4E�RE��em���0�VnK��ػ�s��=��S�ӛp'A���Qt�㭨��jِĘ�����;��_F�j,���C��{���;����N��^���^��
|�w��x���V0b��A=Ekձ%c�L�b��`�%318�����@m����i�B�%{�ZZ'ڠ�����̟��6o�����UNN�%s�J�[Z2��.-UӚǡx�P,�.�}��_��S��wA�pX6N䠡 ��$�V�;����q#f�%��n}C����.��ض��u���g���w��bi�jo3 �c����I��("�/@��s������6�^ŭ��8�"/eo�g6>Aa�7 ��ir ۃJ@� �d��_2J^_��]\h��v5���9}�	�{+D8y0��v��+k��YO�8@׾�ӾJ4	�u�&�I1~{����-��s ��y�U��C��\��@�T�J����3Ȏ����^��yE���L ��lP;�8���{�i��18��Ih��\�_y����DC��`c�7��<�����[��@G�򖊜2= vZ�N{�4���E#>�O�#�va	�ܜ��]�Ki�=+c�/����w���ވ��G�'�7[��
�{C���t�/��E\@>Ń&{yw/��j|�W�xL���ϴ�e���ǨY�P[;����Q�Lu8��A�C��/�Z�E��y.�,]��ea����Y�2n���Z��хU��/�Cn+���'��8e��m�A��3�F����IB����y�6�x3`� �;8SHw#���Y��Ǌ��� ��ʢ��<b$�At��2�K�!� ��D��OȥNt aNP?_~��qj;���d���Ťn�V�ex�A�Ņm��S�����j�s[��橚�� � ��n��=Vs�ws��Ǚ���$Z�K\^�[w����R�K5w����˼;a�vc�3zS�8�룺r�wZ]Q�A	�	���Os�L����U�q5�3i�h5��Ldx����G�ֺN.5���+�����ݠ  Z�Ƕ�ܷ@��SaS��ٸ���O_5��x�@�(s̻z������43�Z9J���+y�u�rBڻv>�/8�VDx�Iz僜�i0�r4��l_�c��0���WTV6�u}�H�R̪�wĿ���9<�����W����,�`$��'RI���1}p[h�UǙD�lg52U�JdMud98�t�	}�DQť�����ag�6Y'�+���P��d=��\��&����w�jp�=8��ź*?`���:v������t~go3=������=#��4>�mI-g��ӓ������>"·Ԇb�X>]��z�O[ ��!�M�f�"�����'��KX�I��u%U�'?=������V�t����d�
��ހ�a�~�����(���\`��l����IC
m./��ס��3>>��}�~����x�?5�.��S��8߉��8D�J�]�[��0"����/j�P�֟�돊����W���Z�TXi��Hs�w´�N�_����;u	�	��LLL�������
a�AT�/??�*���B��
�w������_D)2[��]Bf��>h3�ե�r�Ԣ�E����V���um�Qψ�vS��U]��i�KC�y&�5�� qͫ��" '�q{��@��o?+�Y	����8����#�'٦�ǲ�4�ػ����^/����.����3l|1��@�!�~����n޲�� R$�f���?c�}R��5�;�Yis�8e�݄M--� X�ˠ����6�>6��5�P�?r���S�<����d��p���N��H�U�Wc+[{b�2��߯�(M�^�Ri:��3KL��R^4�H͒���(�~�9B�aI(p�����wz�!w����4������ [!s��m�_$5M��Ѭ � }��QIĞ(|����g� ��|�p3yp��w������Ҭ�,#�E�dZo3A�ë'��e�֭�������lX姹d*�b�/�ܧ%ˁ=z�����;"I,b���*�����P�{�!��8��b���@���ǲ��w-��6%']�b�(#b�=�V���C0�����w�o6~kѭl��O���k����v��WVj����bU��Ѓ���q&� M�Ծq,,e���.�'��$+��6��CT\�¤�V��l�
m����Րq~[��6%�X~�I���d�/�hx�"�Z�t��{�y�2I����@Mw��J6A��'�����j��Z��p�)��)"��KF�[���;R$���X���ς��*U �&2���8�{��C�ZZ2RY��/߼���9=}lf2�)�r��tn���=G?�^�G������א�8K�2}�Zf��ld���X����"�2������S��wD��ˇ���T��k8�3�����cV�(����y{<p��s8Kj'E�p�e��G���7ԒW�TQ������<!b;���Ō�˩w8J���xv�g�Ծ}���?_L��;��Z��8I�;�bxz�ȥ���I	��	�(���k�)>^X
��6?������蜌jS�Z@��U��@3�!iN8$*��o��-+��\{�p�c�V���y��ț�6c�w�qO�^M��%���r� 1D�J��&3���^��i%<�:~,���"�.M�>�A䲬�|
�>~ȏh���7и3��jҼ�Q��|ںrm�!X�Tӹ�[qY���!�߽�� ��n!m�� ��ht>�'%�F�L������	�����:F������WxŪ*�N�+��D�e��VNn��WD?��M��ʪ��J,�W8v�=��ܓ�2��u��]��>`���6"F�&��l�=�xd�A3.���˚Q\$xd�
F��8x�__���}%L���H����Y�2�f�tq��J��GO(�/��L�$/'��ʞ��z{��v���z2=��wY0��)m�)�P�X����D
��.��?+�b$��~��������p���������K�ȭ��b��#�kh��[w3Z~��-i�-��V��{G&�4C�۱J���j{�*�NE��j_��2�t�V�XT����_���|n4��۞ڼ���Ӆ�w���@
T%e�@8��]��*(�Z��e�yYM��)`��I�r�8����Z��JX%�9���DGl�y짬��[������ʹ}���H-�m����ɷis��{܋�}�U%���}d@e�9��۱��XZ1��2�;���0�og�ķ2E"F��Ix}-�T����F���޳`3�B�֓WM�(�~������m�5}'����_�߱wO0qʓa5�	�nps��枞ׯ^�yq	{�X�|~	�U���J�h��V�f[���sa���w��y����]/���Oe���P3^(n�Ɍ��/�6�`�u����&X��g���)	���`�'�!����v��IMg�$����	�5����O-l�R��U��1��f>�Q�w������V��f���`)���`�&�����v�#�q
����Y1��,z}W�I�.�m�Ky���?l���*2 V�֣Lx#s���@��~5�v�W)DFG�GH��H�_y��L��ޟ�kq�=��p��[[Г��>Z	>�;<`��d��"e��|V,�y�B!Xې!�Q���>l�}ơ����,�l�uܟW��2��� �"��E&ZSb�/�o��V�9}%�Q���S�����Lq�����t�@��1/L�:D,� eߵ��|���YZ��f���|�_��9�����;7���zn�~5jN�0_'�b
5K����i����T{�0b�o��v��@�*TB�,�1��2:��=��hɯ_�x��5��(I��zg	�?�ZS��l�4�j��Z�ɗ��[����d�1�8)f���7��?�R�r>��=ف��3)���������\��W��`���Ad������w��/��w]�/:���għݼu�B{��w6c��Hr���>�*����}��$s�ٗ"��{ϣ�4��@��lFF(�k�Y�D��u�s�\v��fZBl�Sm�wpA=Ϸ���l�g�hOо!��Q������)�����I���*H�������D�i��]�!�хO心��F��p
i�� a�D�W,B����P����2��Q���R��Q�~d~{�e�R�Я�'�ML1���-��z����؝4E�D���(T@J�<v��<f��#��{�kr�mK�e���&��%�4�w�%�"���	�F��M"r�T�gxʸ�?|ѣ�3���Z9���a��.�b�U\��������~J.� 9*g�y��q6��K����U��2��&�G���9biho�����?%���!^Aˇ����^����lu�4�YO`�����O��
x��������ۮ�:󛗟�2�ajR9�ͳ���%�
��SL�������Ir��k"Yc��\���`6~����κ�U	�,4�ʆ�c���s����d_���M��|�����X��/�J���բD�y�7���۸ﴩ���أ�Lux��������x�2��l�j{^������(<��R�@M{�a�QR�/z����l~�|�6�����>D�	Nb@JO��r�ui����S��Ə�P������<�&��oL0���I0}���>{�U���K��31�_@�3ʓ�v��-I�%�#6+���&�U��j���a��/��\�*���J����m��\t��T&��㏱pL�vrc;�Y;���#�c�2Sm���o ض�K�����a���"v`=�=p�7���� 8+~~�z=��V�А�a63P�yM�sq(��ny�Z�����=;i��[�?�����Q���h3����q���Y���y��$l�֔��_��L�.�D��M� 15�ڽ���bd�ǿI(�^�#�����\u�e]9xr�0j�3��LG�Qb^�
ݤ�dt�ʞ=(������&O@�==�߳�`e��?u�mߛ��~�iCL�}A݆!��҂�Q��	*$êߵ_LX��4��6r���Ծj�����H��o
�խ��6! �*#� �N�5%WM ��	�
���_w�/ہ���f.'G��|ZBhj���������P��x����{�ygۤY��{�G��he��Pr�^�	AKK�q/�*x��I��^++㶟f���H�;�Z��f笭���_���Q6�����3D�'�8�KR��X�4ʛy�CNi�wEE	�(�x��>ʅW�����t� ]q�]�JR�ۺ�"��qk���-���f�<�dg�j���?����4˗�R�n�?UA}{W�p����(��o�����?��F|+`DRs~�o�X���;=��k��+�?M|a�DGVf$^�\�`�=��0,�%l wQ��b���Qr��-[h,�!�����������-I9@~�­<'��\��xț��ar������"��G`[�W~)GzFF�� �/��qO�^L���_bk��&�
�������H�Fx_��]�i��9	��}ۯ9�c�c�pK��@={�8��K����~��v��qƼ�ֺ�Ož���-|Q�a��~qʭ�6������df~�A��^��mR�rQOՙs���'��x�<�!�f��ID��<]ӯ����tB��nq��Ч88��i���S��$ �2SR(Q�6s�p��u� ���Đ���S����yp;hI��ܩ!��X�U\p�ξb��og����c��l����1�J�8���W�Y�@�Λ������/ځ�Y�b���VdBz��h�,�HX
�B�/����QY��+�=��t�K��tUܟ��&^i�ݣ�j�.{�T��b7�	�}����O���N-,v�z^��u���u6���:z�ôs�����A&�ǆw�%�YIqV��=.0���(�� g��|�����a��foCO
=X2C�5ɚ�2�YP����(�Vh�/��$���!�!G+�1@(C���9oX�n��:ID)Iæ���X�D=�m|\�����s0�2|Z�� w���J�p�a����� �(:..._�k���̓�j�]e���W��Nt�t�p�P��?�����Bi�S^�0�Fr�d�y<p���a���Zn�X�*,J�����ʕ�T��?�O���y��1��+Iw�j�ņ���?��>�եd����WUou|�ۓ?��p����)�!�l��1N��o�\��)1�m�M=�±���ò�4�����Gp�\�@a
�i-��|���PxӨ�c˴x�O���-�-�7�^=5%~.���	/�QW�M}���	i	�����ZD�缆
-e%�C�m2C�ƺ���6]
�<_�J��ň��oU��@�b ����ye�G#/����mP���E:bø��L��S�x�1�e��is2A�s�U���C�@	j�vɺ�xu ��1T�E�E�5�����$����$(5A�؅����������������p5M����,ȏ۪^8��h:q�:Y��&� ����b*�{��Sw��xCju�xC� 8�N�=����SO��������1p�S���,��G��6~J��V�k>m���&9���ZTbF�2�2�V%miQ䖼����Z	}�x4i-�����I���8W�3�&���U��z$Qh�7�����TY��n�Q�"��<��Yl�A��G��M�l��_m
o~� ��&������<�4�����	U[]�G�_$g|E\���EܚF����*6c#%�)o~��f��a���l�7Aԋ҆������r������̗�@�=�Ç>qj�+I���M1YK���W#ÉG��
��m�&k,�9n�9����5��v��X��"R^hԷ�v|y)���:�>+�R����A��=��������y���z���J�y.�����0Q~$�s�����>L�F/`�!���l�E2���ѺJ�JEӌ�Cǩe�����D��$8:�����͘]Kz0~�)��Ŭ��?�����u=��CW2�ه��G7���Gϰ6�/�o>��]��j��%��j5��F�M����]�.��$�u֠��c�����K����j�7�2#'٢���LIK?��g���.��@�ՒZ���c�5�G�HV�J't��ilF4i��� �5�����S^B'�D��/Bìv����'� ,���m&��m�C7�9mgy�X �S�Qh�p|���v���쬫G-���X5Ҝ�5G���$��2���D�l����}���)$�Ȳ�Y�\;�(�p:��(�I�zx�;d���<N>ȋ�j\}�_<}�z����kQl�8e{eu���!��5�$�׻E�9A�D�����j�^λ$��O-�t�܅<x��˜y�~���R��[\c#��abܧ���+42���J��/$��f��<P4�e���\�8ON?j��S�3*����5׳���z�˲�kNpCQCC�Wlu�@�/Er�U�p�l�lAf��SEd�o��f�q}<����H&ِ�Y�6��~i����mg����	-:_w})I���dH1i|].>'��h�L~<�x�J��� ��UBv�.���z�1J��q��]t4N��q����v��'�q�ol<�Ȕ�@�v����^s�<Ӫ�KM��-��2@t���[8/n���H`鄑8j%�З����(��]��P̖d��ِ$1��U3[M�"���<�R�"Dr��}��I�u��]:���\1��%���1���sP�Z���� -ʘ�Hw_̼�tZ��|�Wj57� ������ ��M5%�BP��s�M+��&΀�)����V�S���=��a�R�{`i)�ŝ��-:^O'�u��?�[WGfhh�4(�ؘ�4�ǣ1��{�e��W�Ѵ�&c�Ke�i�D��'���Wa?��_�(`9IczȾ�V��1)�L\�B!���*snQ��>h��a�]cJRkE�Pي�D?�˦�ٙ�VQ��>=L��7�W[���9���!6Wz���'�Z�wM(�j�7s�MٕRY0��6|:9p�Y|��O%?n���Jg���i>��<���zB/Y��J%�,�缁;r�9�y%[=;��~���῍:��5���I�|����A@��p�����AnP�<�R5(���͓�G��.\S�y�H�f@�����L9I��8;94�$��ˁ�Vz|y��r������v�	��=�L?�cυ� �Fi˨���^x34j^@�o��!�G�j�	E��Ȣ,��*VV�N��z���q9'�(DL*��v'X�CJ�T��G��SW���Ō���U���+6Y����[7K��>���k�iT� S��t{9\�����^�r��r�0"Q�!����ͧ�$l.��3�E��k���	/t�2��"���a���d�`z����mL��(�{gW��~�l$����>Zխs�U,���(�5MQ��g��wy�q�E)������F��Mt��U��|����I\پE
�	L����N�zB�{��n������C�c�M.;����/S;;<p��1)|6<��%:py48F961�FL�~]8j3��փqW˪`�|NTggKv�T�2^=�8=����������Z���i%$�c���G��v=�zihq	;�k� hs��ݚWE�S��5����\?>v�q�҆�����J�*��(�"��������C��3u���|���!�/)�5�q	��[��VJwf�s1�1�,��d~��Y
پI`��2�_M�Z7���!7m��V;��%�F�m/�G�0{����L[��@���{��;ѕ�3��̵+7����vA'8��'ײ��>����4�� }V�RC"gjH%~��[c!�nX�xρ���q��B�3�n����̺�ϐ
��;�n�i�1�E\�����I�ͧ֑��@l��^��	����L�I��88�[V��l�r�]�BZ�.�*C�h��gK�6Yn��,:���O��=���l��\<F5�)�=�g� s�����3:8}6O=���N��?&՗�����*,Ϳ�lӪ&��I�Ƽ!��|ꑒ�W���I�*J94OS���.d�R�5m��{Lo�;�h��X�,#)M*i�i��F�頛A�F������Xl},ON��l⭁��Ėo�z�a,0�1��/m\�����<]��6i���.���}��d��.F�&팸:�\���*	J<�-��7��D}�R���$)�A6�FM���u%����Ew��.��+��eO�:�&�V�OjQ���=O~���9n�Y1A�x�R��/2�l���ُJ�Fڝ���$Ɲ�;��;�g���A!���q.
E=�A\Ҕ��(�mp������٘�m嚻���4�_ȥf�/F�jx+�����\�졿�nа�����6���C�#�<���v�ZX��ɯ���U���l����D#�g����i`I[f^ףl�=%�Ɍ2a�_k%�ӫc��ݬ�mY܅'=����߼T)ר�0���9�yg�����%/9����%d��*���7�no��/jrVA}4������V�e;lHu�����1L%z���$��E%ߝ,5�bU��[�T ����c�~%���-c�c=Q"��8):��ğ?u3��AA�f���⦿Y��9��Z�Nt��5�|��8/��
CJJJ�'�7$Ǯ��E?��ywV0�e1I;+�I	��V�^����{�5<���Qy���a�=�Fd/��o��Vv���|�1��xo𔺯P��Q���L����y+D]^��-��^��S���V��k�:̅��ւ���l�`{k�h"�T��@> @�UP�XW����G{:���#�3WG�Y���{p8O��K��?�+�W�R5̻��;�X��-�X��_���Z�i*���ݝ����jqn%���	('.��M��2���FC��FÐ�u.���rt9��ye"W�:p�
�UP��~w��Ck����VB
_Ϧ߅�
?�B�m�eQ�0R4���r�,_���@2��S����}G5\לM�1>F����6����X��6ʁ��V�w'�M���z_�n���i7������n���Sb�����n�Ut�jX��1F;���b�����|��n��]�s���&�)U��piƬ�����YB����k~�����<υ"�L�����ԇc:�}#-�d6ߴ����fv�h���ܹ�Ff�P�HǑy�v=��S���h[��3uR*-�����i�J��5r�J�}D'�	���d/u/�j����(��v���3dد�ã��˓�[�*u'^���2,���A@J����	����$��n��e���A������������.x�㬵�>k��z~��yI	��C�iD�RY$�bu��ܜ/"�/����Z��e�o�қ�lM>l^i�,�ޫI>�ն�+�ǭ�����������6�j��o<=?����\���dp^��쑖Ο��]]�0���T�z"D���|pP�����5�^��{w㔜�6�@��8_T��
�����=<��p�f/����u��;�U�Cv�l��\3:cxؘ&�B�;��͑��������na9ws�qG���J��bٛ�e��n�0/�(�dqG��H�`iǐK�n�����p��Y�I�L�XV�2�}�0x�Nm<�.rx�O;G��;�j�!"!�k+�~݂�0��xU"Y�E3�kx��81���ȃɹ,"
m톶B�1���C��s]�j�|,dh([��<�:�7QV�CQ�k��+g�$O'�.*jy�]�1�t�1	�_x��߇p��y5�[�Հ{G��z���|7�oC���!�4����C�H,�a�kļ�V��3[*��J��~��3a&�����7s3��
w���җf[�!��YL��kD����ܛW����i)�!0�r��is\pMNE���gjP�ýV�7�}�U�|�]��j��&�m�˰`��u�X�ڱ�G>Rz+�Fc'8ϊ�:s+ۛ<�8p�9A��ڛ(���Af��畾CeY�zw� 0F^�4|�N�{�y�T*qlr�%{�V�q)�:�(=����yzg�F�G��kJ�P��K�>�v�4Xd��e`}6X�Ou�7��g���7�VĄ�����&=�7�����K����<!�'5�a��¤���o ,]�����C���3s#���7�{i*���� b���[b���o���hW��PZ��_G\#&�̺��_�/���mh�6�k�}�	�7g���`x!Т2�Hj��!��൤��m��+^O ��E��$�y@@@���F��y�ݟ�rQ>�hiko��Nԉ"��<�����R������0[�;0t:�����ygR�,��W)J�rka�?�lq���+��������T��"9����o���xB��j�sG����ׇWs��U�4���HJ&��E���:�E����w3�#�c�YK-d9j1�S|��[g�J�w�֏�t��!S&�.H{5�'(�"�r=��D���!��4po���͇�=�]�q��13�aA\��.�;�����>�'�e�k뙧�� ��uE['���7
B�X�"Ja�3�1b�pfWB�p��p����Aw��rS�k"�˽�$��r��;^�Bu�2��h��f�D��ui��~��C�B�YI�i��@
# /Evx��Z߰WlӪ��=X&|���d |4���9�$U���W�Zi�����I��y|� ����pv��,�0h8�n�.��n<d)ȿ�����yJ@J�)Db��lw����o{˪tX�8\|��C������4A\c�����Dm%H�Û��%�y�*�<ǌ�<*`�K&�~��y���L���Q���j�����|*iG�<��H��E"%8�����C���	�	��G[y�V��C�����,P����4�O#~C^�(�7��h�q���Z���a�I�)�(������c����ɼ�ɨ��-�W��pW����ڊ�_g��2r���|�� �*[�����7f�c��Y2��e����If�c���T�-�;
ƛf{2���/��2�-���yuY<,�Y՘�1B�3,��y+`�	�e������;/�xx�N3ws���h��B�,i��c�\�;;�&! ᇱ{�GS����[�j|u�Gǚk�};�ܦ�<O�
�F���=vRh�)��M��ᱚX�kҟc��PжR�CKn�2θ/�Q@#}n��23�[�G���A��68��b��L_����Ӫ��d-5�A�2�	�Tϵ߿��ՖK>V~LđQJ����<9�*{�^��|_]UQQ�%�� �0���Y��'{)������Op:�����<�����ú��y±��)�W;��Î_#Tn�:Z��t�
Uh�I��"+������j��$LZ���\j��� ����	��?Ə�9�kMn_�P�+k�^<�r,M�]�_@PoB��qR�DA�b<�`*Lb&|?00�<H�^?H����k���h�:\9�k�e�����z����p���M�Q�����v�ͥ����Oz�K�ٺ��m�׆o� c�$�AdS'��qӰ�&��X:,�o�A�IfM�F�-������%�,�S�!�`����0T�T�Y��D(���'�!��S��ي�)y+�gA��ݖ����hH!�ċ����Ra��h����$P�?C~���Z	DX)w" %��N�*��H<3n�A��11nƑ��k9��[P0��$Μ����#I�]vHcӳ��a�����X���E���<����9 K�U��I���r!ޔH��n�4�+S@��7^?�q� �6L����3��p��ǌ�q��aG���F=a�r߲��2]ei�ql�1s�	����v�>��"���s#� � �,�YYs���������dU"�Wo[���WRq�L%$n�6��xt2��$%#no�`N�yq�!<�Z&z�6A,���jc���
�%��+crAf��V'�͢^j<�e=��_���P�Ǵ�B:���d���?��o"1�/q��q��ҹb��kJ���{$V��ͫ(z����'O�J�M�[��*'4Ī�� ��� Q�BlT�i�5���Ս4C���+��a�>�k�"���S�P��ZւQ�j���Q��y{"�����w	�B���n������SOS�(SJXE?��iy3r3���3�a8���?NQ(�ԝ(�YW���������"x㹡�Y��G;[�F�y�~$Q�4�5[<��^����'�������ٽ��S���x�S�����K}���X�����܁�N�;\��:��a�#����<-M��,�E�^���^��Z0T�����= ��ZZ�����֘rYE�cȨ����&������@4����������;� �p]���oL�6�8�q4�414"��\y�<6k��yjzm���Jy�~6��C[��B��~�8����ʸ���{�:o$�1~��k���®�D2�����!jV)��Z;�KNX��Vȼ��x+��V�)���� ���,� >���뵄�����(!�� |��u���%��?����^��¸�6��P �ڋ)4Ԭ������)zªG>JL�SR{\{V�2+�~,)9�65��{��W �lEUU��"Τ�椮wt���H���Ep�cZ����z���f�o�+�O�9�\+�ΎEI}�>O�'�e*�ij��Q�P��Km�� KZf'5�ہ�'���π�/z]-�4R`	m��뛟e�b>�'��a��|$�u{�X/m��,A>�z>���f�<ޟ|���{;tN� 	����Jf�ۤ��UV�,�窫���<� �NkV��I �5�E��,Ņ����x*YR�2`vG�����me��k���0��~ٛ����-�S�f7K:5o��[�:��>8���p#K��\���~k�L��\w�1��
�����4��$�|q��D�S��2���m�o�TaNE%k��]�eҀc+�o/*�]#sSѣ��tF�WO��<�&��b�>�av}���<��R��E�T����q4b�;<P�ԉY���97K]p�e�o�_s-T�c	�}��%��b��8����,j����z\�?<�?�����y ���sv�"�b���;�8���;5Z���a�w*�f0���"#/��8
�A�'�
	�{���4
�������-:��I���d�(��M�]�ɦ]h�Q��-S8~u�(���ʓ��Y[����Z�L�"o���I��w���ʾ.`ބ_c�>Q���L6��!�c�B��+��3Ǳe�d��w�4��Z�Z?'�3[�Ωab�j�zQ˄��d����>�gK�43ߥ�~n����d��OLrk�(��ȫ��I��ׇ�?�"������y��x	�;��۵tXt���f���$<�D$|��s(�f����v�roez���)z���Sv^�败�ʗpv��=���+�%��ǭ�h�KLu��c������� Gw���YB��|*
��N�ҍ������q˻�S�M��n�dٜ;0�P���;�:o��9��<��*�Zy�:<��?�1����H�Y����mM'w�����2R�D{�u#����\������B��n�w)�zY�/bu�3_�Uy79'�{ﶪ���Rc���������[Φ8rb�$���'W�~����P��q.*R�����c�ڳ�G����Z��2h#Y�����=��T+�Õ(=a��kzrA#	\�@!�z�[|�^�60��~��a�f�"hL��R��o�����>VTT(f�	�J�m�B��yr�/�\w���i���G c��nC׈���ν�M���B{��X��ޯM}j\2S����ٿ��_�kcd�:��g��ml���S����T���qS*G�v*Q�j���]�q��uY�;u A? �O6kDA�j��ﾉ�d���q�A7�<�ڜ�Ja�����V�i�Y�Z�:�]��+�S:��Ӊ5U��S�B��q[l�Ta~���B�S��_�n����|��5cK����j ���f/  �5���3ı��;W��ؘF攽��_������YX�d��"�˸.g^��n����ŋ�{����{F����xi|�Ъ��m79ظbXo��V#W�����1^�=x�ΰ�N���O?uu�C �2&-��1�i�c�c��Ăoo7����!UUU�Qr~-�_)9����s|�"zᣅ�
f~g1&r\D��_��ߥ�w���GC�'02�iǽ�^��K�ra��Ҏ7+q"W}�m*�@D_DF`_�S �si�J��R%���Ɖ}�,��e��u�n^�G/�åN��d7Oם	r4�tq�}�j�M��­�0��-�I�����7lQ5�u���D��lGD��2�p_�0r�Kԯ�+��f�Q�e9�v�-œ	m�6��B�����/��q����ty�\d�Qo���D�r���s�$��ڔ��@���6	~������Oh�Wh4�(��0С��}'31L�깋�����[3�,ֽ׷�O��Sb��
�m-��B���O�||����g�2tL0b&j������f:ݲ�۲�o������o�"G?
ƅ_T� �_^!�P�h���S���>������ήO�Ϩܡ!.\�2|�+��(�����46�k�⦻���l�vG�VF��0ț��gu1�^��0%BR��W<ؿ6�ݢ!��OM��L���J�)΀�.V���������A�'�� 9� ʇu��!��\Z�Z�'N�.�$p�遧��Mmq��}��U��"��i�֜_2�6�ܓ�x�,���C��?���U���������V��Y�2�K<��NM ?���.\g���7��R�Q��v��h��呭���Z$ֿ����un��[W���@��T�q�|���-��=k)�C*�|���")�G��Y���9�3n��z�$x���D�o�\�]e��fQ\L�g.�}���(�������k6A��R�ǝ� ��ϭ�$���hVu�&��V�#�	��A=yh��`�C�/а�����o&��-�!��b2�Ȱd�x�.!hJ���o�ı~���nL�hg����sQ���O�k)�j���>\�b�lki
+K�٫~L/��2T���=��Ǘ2����ug�Х��6-q�� go^��A��@/����q�9�2_���f�Ӳ�� �ji��u��v3�=���J���Np�����-c6�K3�_t����R��-�c�����7FU���Eh��K:��G4זS,F����DE:�a�3a�#74��}�b&qR�N82�š ����?D�wR�&g��-;;C���p�e�h�2vgg�V�"l�>Ss���s�S�r�y�K� ��:B�����R�ps�Z������!��_ݽQmQ*����u�����Qoc�J�e"�(k�d%���r�����Z[[3x�������r4쮞��D��S���I<[�e�d�1���������SD1l�LΌ}�
�|c�d��˗��Zz����	?�r�<׸�/o^��c�r�F���f@`�Bg�$*�[>#e{�,��"��U��Q�#�5��"�5Z@˓ �`�k㘽%�NБą�cS��N��[��4��|����>X\{7�D;%��8W4?������/���B@�psC�A}��7�������"�N����_I"x�yP�>��!1�������ڻ}JN�؟�ڐo:S#�u<�ӈ�h�ϵvv;�L}�Bծ�66B���k�4P$~�E+zM����9�2�f���pX�CW���V���q�����gX�����NEnw����90^��1�2P-�x����Q�8H��ژ):������bǉ��;sw�^"a��ʨ�Xm���-ʳ~� �GB���.���d/�)|��I��w�}h�gr�g�KF��;��=��t�v��ţ4�W����DI�B��,jN��B��Y��Lmv���kd�=�W��T<C"���/���@�# -�y8���1su���t7R�8�+�����{W������,�,��H'�:ﷻ��w.\��m%�a�T����g��n��1{�f�{I��v�7�^���}^�z|*& �t$����hko�;����bἎ�����Z^�c�,������f�'��� �*�7,�d��)�!��$�@b�j�hp��L{�#Xkldw3���$�..^W�C��L��e�S4�h���	�����{�>4�gS|�SN�M�{W�ۯ�[z,�[��8M�a���>���2�si��F��.v���T�5����$V�k��a�G�=[���͍��B���V����V!G�W�؛��e�a|�!�X6!l�����}�"���!�hgWU�M��L�-:��F���>�0���t�2��~ReEA��|��C�w������:��!+�qރ]6Q���Jn-:�2:�1��xa����5xm�R�R���_�/ϕ����St��W.��G���֭r�_�quD��u���`)/�A�����ۘa)�I���������i<��q���
��e>i��rvs]�P񥺷L���(�:����3��B.�������T��ܒ�	������0�����`�~�˼�S4dG�5�!��f�b�{��ƈi�r�?B�ܳ��6_����4�{r��;,.r�sw�I�K=OѦCb��E$(�&�GT�Æ+n!�dF%'�ߋ6�L�<���gӬ�ޟPUR����򰯷^�G��I��1�<���a�X��>$g����rww�o'����SV��½nlM�~I��_�5*&��9m'�{��C��|~#I4V�'P|�J�G�'Bū*�&'��͞�ݱ�,����%��G--�Uv��PL�~B���a%�&�� �,A �h�EԷ���h_g�MKT�ط�:������`)����Q��l�b�k��HdT�+1@|��~��"��c�}(�S5�����ڷ��>�n�\�7�� �HI�G��{���ú�SJ�'u���gJ�.а�����VZs�Ke�)�/�S�x�_�s�ׯ�~��c�pcL�ٺ�\�:���!��%�ʋQ�@ޯ(+�����V�<�����V���f#����귡Ǹ�l�nlX�l��lᴗ�Ƿ��BB�����{"X_��X�T/'����Q��DW) �O@��H�4�^�0`�h 
�^Gou�P�6�߾�@�9f�[ў��(Híp�&���xt2�b�>Nrņ�`�������m�k+"`h:�g��{����)^��w���w:
^B��?�0�M��K��0M���r����z#�)���ڢ
�z����c7@*a(�� ��K�A!Jȴ��x�W��w��M�}�ABѻKP�C�r�������*�{���5Ӂ�J������ی���"V��;?6^^.�$��;vgz��X�/I ƣ� ����Ԑ�f��q7|�|jRy.P��}[�{/r���(�p�];�ܓ6$�	q"gK3,<T�0����7�;0m�u��_�
�ȇ/",����N�l0�0:k����;q\Ee;��1cotɩ�L'���[��.I�8o��j�݀���#��� �h��i��@-���y�>K�}g�D}��Yʟ>\LZ��"��/�;T��ϊ.ERC��&r�M�-Z����O\���uAc�c��:�U�fNО �jɔ�W�P�~7��������++� {��gS�ѥ��s'S�hX7q�s�ѷc6D߲��(�뭇��A�Q`*�Ok^����.�����!O��2b����<�)��U��X��#����|��|��e�@k�C���ڏW�C��X�/���ΎM����`f'BB{{�Gg��]at��qk�.؉}��~pX��q�s��B�] M&��Zo��;B�[0�Z�\;�nDo�#���E4��T�Z!� zS5� (W����ݽ1�{s�
p������_���yQ���;�1Ҫ�fqM��3|��+y��c�fs������NMc&;On��_	B>��sc7�T�VJ/�5����zD��f[yw/I�����9dd}S]/1^�t��8������g��6?�1���8�b�?�2�Fp�l�V�$*JI?��SW>�@ݶ1^��~O���q~c�Px ��ʲR&HT�GN����vbS�8~�^��qBH�qr3Il�B(��"���޲��u�w#���mO�E�P��� �å)P ����׃�?VgR/�j����d��`�/����Fr.cC�3�d�V��~��}���/�8��=P��g�qQ��k`f���<�Fw�1@.������m���  �<��'y;#��k��.�L�����U̵�UضC�t�v�_/�j�XTG+�c���^4���ͮ8-��o�� ��ST�y7(i��̇r!�R ;A@�E$���w��W[)��^����9�f��Þc�,,~�߬G)�>h�yO����A���-+��D	ģC9�l�9��!���/�V�I�vq⦩��$ߥ_�ŕ�fT�-�R֔iJJ���M-lP�@�AF�M/IU�[/����ҡ����M4x�\U�x:_�&c��6�+	���VX-��<�厅A�����ֳm|&L}4h���0����ȿ�7@����.�~�0z��ɸ�-��}�#��S�k!D���U�A�G�^��$D{_���W���<Xm�=d_����YsYQHdx����v�&�<���1mX3�=r�'ԍ�������@��@�=,O�����`��l��&[��7��\�����+�����M��X��k������W#���ND�{��O��P����7&DO���p9�������M�"���$Cy�o�m�Rubw*�f����O�Rn����z�nY�-���&w9�A�3�r��_�<�gf��Ty�"�=n!�N�Q=��d�:2�����5[��9I���Z�&����h� į6�s�M�:`!v��� ��{Yr|v�#'�pq}�E
7��3�z��tE���^x	�L2�~�,���k��Z3Q�(�����->�,[�0���,��Ib�׭jq��yvb�,��
�rkX�r�x#���z���e�jKɉ��l>)Qd$��~�]�rp�	dd}�s4d#�Oe��`)A�@'��t��B%K��d��������,N���e����%��ϴ�O3(�~��Bm��ײ[������ʏ���5Y�x�J��=�9<��sk�h�9�)Sx5�7{�C�9�]�ő 'NS��O.�g�/Ц~F��i�2��%���Upv^C� ;���a�k�
��6C[����}���od^|=��m)_-G�[���ԍ��Y��� �7~Y�vNտ�mՀ��X���cW����
�L���Y����FR1���b��b�q+C�?k>�$q�������4��si�E'��g�t�q�:*��8/��vYEMU_ki]a19��6�JW�b0:���b��w�S����;�!٪�9�ا�$C��Y��1P��L
�� �fd�VI��7^!�t`pc���!�jf*������WjOS�7��|7���ķu��2�� }����qMg% 9���4BZ�
������+~SD������k51D�4��W���&Uo�Z�K�;U��4�^_�C��=%I�]���9��5�OO �N�X�A����y�y�[�=�B��E�'�|5���J����O�u
uN��l]\��Y�p�܆�~)�W���C����;g�?�d����Ӥ��o�1�����qۏM��ͣ!�mϵ?ݢ�c�e���յ
HT"��*�B���Q���FJ-�ӵ1�N��#��� fc�?�(�9��ΐ��2Z� �,αςxˍ���2̽E�|�0 ��D��`�1j�Z�y���Į���=O`�seU��ҫ�:`�O�^SZP� ��Ce~�W쵹��`���M�����M���\o	^�'u��#M��p��ó�%�?��W���3^�SL��~���Ϋza$�d��zv�ʪ�X��^g�*/��$� kv�#s��"{����Jѻ���I�Wº1�3�d����x�U�w��*.|��Bճ�����	��e�7"��G��q��wK��b^�y�g�1^9r3r�?����QϿ7���N���R��Ԕh(2w�\+�Μ�l>�OI��a�wY�?U�;�R4ZΝw����ү�;����^w~��j����ZS!5�;�k���Ǣ���&.�6�P6�+�
|���:ZY�w��&��zج����MT�mrn��Y����?7M����E�M�/��~K"~X��8�"mx������k*g��~�~+�����^*m�#��,�pc3x�抓?��\��(KC:2L�\�"ٗ�&	�x��_��'�5�͈�_�ըB�㊘l�W�wg�BܰI(����Z���t�;��I��~�W.�Jb r`���JQ��H��^#�����A�ǻ����%\�'ܾ�,��b�6U.��uD�ǝ�g,!�G:ӓ�/���.��se/11Zǃ�1Tw�F~uPy:��H��9�;m�{#�����w��cc���(�je9�����Ɋ(�~{bh��1�3,1�(�N��d�JV�#伎;��i��@�
��M��c�`9���8�ٌ�*�.m�}���I��*��P�~��q2gex����l���������C�\�!��x� Xp�� E�Sp����q�����Z9���&�hW�_7�.&.���`揁��&�/%,^|��"���Ûw8��!�Dԭ�Ж��Ϣ �f��:��w��/�Y�
0��>�%���@�F�W��|w0Sto��bd����U�Qb�������N���F{B�����4D�6�"�੶�ٓ�"�W�Z�m���b�޸�v挿��w�����E9@�n��9�͔�A[8
r��&��fdl��I�Z��Z�5�Z��jj��*{�ε��am�^��H<*�Ύ[-NT�F}]U#;���2� C����(�]�z�@�W�[��MPT$�9��1��
s��1�i����?���w�� �J^��Օ��9��۔�:����%�2���C��F�d~=����QF�FE'- ҉�2��&nw3(�����P,Ρ'��Z�v��%���/�F:!3�B���]^���l� -�002H)
�Fs�IՁ7�6���AA��ͥt�M&�z��g�L¶$�����σ��Y�m�I��%?�t�ߕ�זFG���'����Z1s�
Q׈s��Ÿz�n��+"�W�E*�uSN�1���S�>���X���gѬ2���_��=Y��τe"�W�����G�p�Y��]�����I)Nr�:S�(g'�7����I��v����)���y��E����nN�pZ��?�D)���kخ��p4:���TZ�'!�3)^s
���z�(��H�$;������4ڊ;mȁaͥDR3��a�\����yU�=4�	�_�;��I���EUb�����ԏ������#��p3�0ȹ��0��������O#-֠��`	V_Ԅ@Ehv =6�:�f��p�9W�ܑә���o�s���G"��ɨ[�_V�^�3���q�^ܜ���ZZ�RWzzB:o=���o��3��=��s�6r&[��	_J���vu%�_�!���x)3��,����Ah��J܊�L�)-��+�p���'�}i�:� ~��0Qd0u��<SK�_�Z��SA�[.������[�"y/K�����̷ii#�vӐ�e"V��U�!j�b�)���2]��~��=K�tE�����U_Nܗ����o ��_L"�jUkV�)����P�D1����=�_�	��$��Rm���<X[[���ʔ��9��'\�z���S����z|+CU�S�o~iS3��ia�O�p��V^��B��x]�(����)��ʏP���z�q��[���+�}D5#�v������Y�T;�K0��-'�2�l+��̻!P%)�oDP�{B��҂i���ɗ�"?Z*I����ň�u����E��:�-�@��C	�H�:�,���D�1��s%�y�l0�|��o��<�%����9w�y�B��I{z����J�o�[�<hg���"|Cq��Zr�f��~ZQ��� $�nĮ�� �m�������[$�MEQ�^��6?�}�o�I�aW�۰<T�`Q�ݭ����M�L��p�2����ͬ�	-ނ[7UQ�v�-��\nߔ;�5�W��a��`a�8�PL0���y���ֳb�5"3���(=崋uc��`qL�*�	Οͺl�p�Q�6*�́�lqq9)��JE�y���ZX�0
 =�xB�:$�ĝ�xyy8㰙/..�/&D��Ue��nS�{��O�Ue�/m
ѾW��ͳv0\�\d��?�4A&�^�k�9l���g��I�y�3φ�����CT,,,%�U�ԕ�n�>JV0�ݳ�n���e:�Eʽ�=���0X�_�f}��g�yߖ{9ݎ<v�]<�����Ł6�0ʌ��7v�W��Ύ
�㙆�+���F�@ddwǦ������tj����%�!ؗ����e�,�ɓ�W+�{��lx���ht/��J��~8�	�_�ۜ��60���{�2?n>q�7�w�wR>��D���?}�|D`�?o:�=����{A���9�t�յ�h����"�;9�%D4ז����Yu�?S|\2Y�Ũ]��y�ͻ�*1ۂ&)9������[��h��]��|9hf߱v�Mf�8�[����l�Լ2G��S�P���NEe�j���׀KVl�x�`i�#O�@ET�;-���L�f��֛2���3����l�B���v�m�_�	����y�'��o��}��P���&�Awy����qj~���M��������m�{�����׳G|{.|+Z��j�4��ןx��>\�Fx��A,:�#���>e��v"��n�FvW�ju)*��K��& ���`��S�k���zy���$Ņ��ԕ���ӱ��k��=!�h--~2x2�Z5'h����V�kgGO�|�M �t���X�d�,��Tu�����9+N�����c���,�����h��g�2�i�`	sc-�N}���\��=xk-bo��BY����*�M۵�j�uN �]y���o�В��L�����-�i�]U�/�`.�}K��gR�\�Yk���7_�����k�Zy2�X���04��.`o1��ϭ��.�.V�t㵌W�hQ���8\S,QA�*n�3�.�)���b�+`��Y`��A���~�ҫ�G���Q��ˋH�ڧ��Nf��\pw�v�őd]Մ&Z�Uqd�^'����t�^7��¼mg�q�������������ü�l���-<�F�/n��&�{�B�Ы����Ij[�����~F�7u�T���a�d��B����`N��4��6���'�oϴ>������A冐�~�<p���w �ͼ���,��zaŹ!#u� Pc��	:��n`�?�,��6]Q��F����^x�Z,׺Y�+�E��/��N+�;4��T��B�X�T �*���􌚨G��UDp�5f�7�|Q;s�<���a������W�$F�q��7�4�@7��" �h���*:�<wa�G���۶�k���=,؂Q�}�WL�hp������a0"���y�߭�r���7A���e:�5��$�~�����*��Z���=�K����(�g^����l����wD>�x�Y��l�6�k]��B�:��α��u�7�<�VF*63Mb���n��B�m�%i��f�BEz��	���� �ls>#X� �.q�Ր�)�ul�kʴH�s���Q�A�&H0��;���=:��m�pQ:�����^?t���޷�N<V�l^�k����EXٺ��;.�o��zYwƝ�0Ư���DK&
.{R�V0������b�ܳ�N�׻�{���b��v�G�Y�B7k����9���/���^�	��ԉ���os�����0����%��Q)�vF�/��wY�&��WlXu3�}8%a����ž,�?��uŹj�*�'lN�.�U�,zKֺ}y�ݵ�?��<(v[IjRc��a�+dY���	h]m f���m�g�^��?���-�Q�uL�yBb��޹���O/�����&#|�V��=�hb�ǡaK�g�ӎ�Cay�p�O��Mg�Zb2�n���}o��69h�����P�S�lFlk�򿾕�8ϯ�8�5W��d��-�<�U�����]t����"���yȨ�^�txx|�?�c��p���Fق���ך�Sކ`�E��:0O�����j<M�u%1)�"S_<P{7�O�\������q%�aI+��<A@�0q�ҧ��W��a1|}���C^z����uB9N2����Y�əq4Y�((�54�>�B��l��l�se8���L�x��+'RZ{�		�Fp-��|��/��?\*y|�A+̅��GQ{����"���'r{%�zX�6��#x�E�c��J.���@�[���
���}0��-7��T�Yj}-A�CNg�NX��샩�%U��X���ȣ���]�[;���x$/F�BP�?-��4������v�����5�y�C�nw�kg7�0� 8\%���	�+Q�W-B*������͙�a��G��ԛ��!���=_M�h|h���lĐ�=T��Z�ج~t��sJ��D.���S�_��:<��E��wO�����uU��0b/3���+�FN*��M@�_��|4��o�����l���2ȱ��\�}�kE��	Z_�k�{;��3ӿ2F���%���Q�C�n�/ևH�!�26�{������Sù�	a��j�w�T����Pi[q����45����i���Ј𝋑Y��2;v��moo/���s	ƖT�E*��r@\^�a��kF���b�K&������{	�o��}��ct��&�g�-��1=f����וUj����y��� ��u�	y�wp �(�/9�\R�������l��ԅ��X��B��k�Z'r�8��Ki)1��e�7��+���ѯ�>vh�����Ha��ϋ���$ߧ�ׁ�K�V���r��Uч���/(~ⴇw��Ŭ�����@0z������w��k_o;�&�<8�i�����?6H.�L�_���򪱴��e���M��?�Wr�S_f��� !K�	���㙁۲�,��,���ѢơL�'����e��Z��0��|�	�(���5�F����-��j
Paܵ����r�^�x��������=�U_�������y���M���ECx_��к�]鉼ԃD�e����o��W ���[�0��Z�I4X�b�WJ���t岱��}�%m5E	/�
��m,�� ��jֺM#tG��������&J�K����� �����ɵ!/uQU+�J�Û��l���S��O�<�I>Y�O��{�छ�<��O����=X�g�7;Sl$s��Zd)z� Ia��ݢ���=ڸreE�~x�Ǝ,��$Ҡ?R��q�}���1��=?�x��6,?
0#�h�lԸ��y��
��R=���8'i�Ǔ	�W�]��7Ҧ�Lr�t�\�|���;3.���1ki�E�F���-��O��J�*O)ahe�G�\-�,�6��51��S�Ŝ���f����9�b��D����ﲔ�~j�=���^��9i��f�~���}�a��K	`���	5!�����-�{��vU�R�*H��M#w��C�i��P�)i��ςDRqh��dm�R�7��'��rOk�����o��,��o�&���3���v�Z6�B"ǔ�F��I�/>S'�����n�a��Z�q�����|��x墅�ؙqx�叠�Rh*�NQm-&���eF���6��z0*�QO��;��[�f�����o�מ
zi|�|����1lƳ���|���[Oi<�4���v�GYd��'��'�:�xc�H���݅��*�^�iS���
��:�h���9$����wdN�Jg���Z�����Bx݃��Lm8�~c��v/<���X��O ��7nUī��\��$��*���ϲL�M���b+�Du������m6�Ҋ\v�^��s#��)�45&,��8�*T0���*N6Q�k�YM4����{T�����h
��\n��pJW=5���4��C����Q�����Pi��$Gǐ�n��nD:��F7��g|�����{;�9��9�:�h<��� ��z2ֽ�����������/��z4�� �&�۲�@�$���D���]4')�0����x�Ym7=�E�
p �.����/��^������8��WSߐQB�,ꛖF�D ������zM��b��/K���;>(W���N��-��������d>1s�R���lIŐ��.9�Zo�	)AHh���h��<�	�c4�TΤ�7�7z�����)>��z���[,�npN��O"�Q���T;l4�<�c���k|���|��Q�[)��QpDI��Gţ��%b�3�y��e@/��������;;g9:�k9�D5XƝ;D��@��5oi���
���^����:�6�r�QZ�܊����L��7 ���V�V�.�&]�{J�s�2$��ʊQ�n��8Q����ߗ��=���F���/%���Zjyw(h�p�PV� tƙ:�p-V��o�� �"t{�k՜��ly���T�n��y '�R���u��!�I��.��d@��hY;������ew��T��ڏ��
��Ga���������{4�I��׊Ȧ�}�(

hi�%�o��N�6q��ݻd��G����2��/�'�^K~�"E��LU�� _j|�X����$�<��K��߻S���6cUa;2�4�#��{~�$�Y�?B6��v�G˅���^h���!����7�&D���"�_qYK�}B�ҟ8Ű��I$Y�z3�W���~�1��4��	�$�M%���e>���8����{Kfw�LR��������ߝ_;��Sk�����'��ӳk'�1WlLQ��l��`"�O��m���RHY\Γ���ۼDZZ�9U�[�Tz��p:WO��ܸ]�<��7]N;?�����GA����x���(������H�y��Sx��nw�S�Ŏۈ�p!�C4I�(��q���Ɵ�	P��.� d�$1����B�����^j3�	��9K	Q��<�=:X��ځ����������.���֪]V�cum�ϋjG����Z-ٮ����Ӷ;�P�PiP�<S6"ȣ��(0J1Sˋ�=.Dpn�譡l�>ja���3��m2�dJnL�[h��G�yӯ0u����x�,H_�ҭ��;����x�);W^
�T:�H��~��%�~�U��.�h��Y���ɍ8�|���%_h�P0��a�Ƹ3��!�Ci��b��ۜ��.1��@�����4�]R*�o��$�H�T����p��*o�x�)��}`7�������㾵��6u����@���j\����d׏C��QZ�n�/VO�ev�t�h�b� �w�I�9����+����:�j�*�Ep@��4��N�	�7RL[�z��x���)��FQ�č�8�|�P��S,D��m��m���q��ɥ���䢞�X[���� @�mB:}��[���y���N.�/���P�����3���'v�qye�����щ%h��V00�Zu���g���_kC�̱���
��{ ��������n�����'��g]�M\[����O7J�CI�nF1;�rQ�U?��9�S�������4q�����^��B��dyy?S���G�t2�:(�	�+�[꘣�+7�FtfgHri��j��]m�[ I)��9>���aJ8�����B�b��@�
$�G*r��L�ˌJ��S����}?�0����sc퀧�ߣt� ["�L8Ե�`c� v�.�H��@6�5��m��v�}�����y&�8�d�}*S�=�7�1+7�2�p��?u�=��V������1����\���P7�RHvo�+I)��~%�|؅�M�%;M�Oqnɬ�}36g��׳�����a��+�ԫQal��a���$b �9ݻ���6�
�3bn��\��:�G}�m,�u��܏)L��bQph9����y��4�
����AR��yR�b�O�\���,���6�իv\�r�=�=y�/N��f$�z�]D۝U����D_�����sZ��E�M����0ϡFg�N�#�����ԏ�[��$��,���1���?*��U%��>���e2��7�����S>�6\n''|�c�l�A��z���w>�x�{6�s�dax#��V	� �����M?��FyQC*1 tb�Պl���h�<6Jz�im�񑟷y��%
��؍q��H֌�����Oٛ�vE)�6��"�\5 G����y�T�1�/9���J�2�!7�}���2��Ä&�qU�΀,��&IdT`�����Q9~�xXZ^'���ީJ��R�25MX,͎��1�:�c��~%�995��°���Li.�F���{���Tp|ݪXc�7�,8b�b�Ѕ�UȤ.�s5�!b0S�� Y�w�<2af���)�HPET9sP�5�7m~(o6�K�@�m�#Bû|*�RIQt�<)�|�Q�:P[�A�3C0�&~й��?�>��͵����U�%��w�f�i����-Q���<�=Be�{�_����:Z�m�*N�{F�����V�&*�/{Ѯp��)��M������ٺ~-g�����[�V�ǿ�� ��ڟ:��w���DU�ǻ�ǗY~b�.vr� ��	915[P��Ɨ۽R�Ao�I_�-�t�sQ��O�*o��������D��16ܶovVôԤ��Qy�%bN�8���y!غ[���ѽ��I�+���.9�_������qE�rA����?3�j<~�3DAe^zڳ��-|�W@�(YR��xu$Ő�"���.�z��[0!/t#lc_��F6
�2���r�~}��t��P_�ZB�r���s>��j?��c��WtD�
 �G��Y��peN��ii)�PA ��&�[�p���T�M�
�Q��^s��}`��H%�d���f|��F�:�ܩO�T�e��ٶm�N�h�.�F���v<��ll�V�k'ӭhDf�Z1P�aZtX�	���ǝX�'Ϣ�KQ�f����0Ƨ�ُX��ߩ��}�w���ƺ��!:�t	"��2�Zw�G�=~X�ܜ��j-��{wQ��Ȇ�"��תj�ܞ��|cm�9�Zz4���!��i����[AIH�Ц&2� dD�n�U�_̪�Irg&�3�H�Q�)f�=��?�L�̟��6��
���ȤDϞ �����8����Pp�N��T�椧w��d,�;B[g�s��#�5���V^�� �K]G����r������#�o�Qj�.y3�N���w�鐹z��S�� aV�R�_���b>�eG��������Ʀ�Zo��D���Z_�Hmb�k�39�[��Uv[�����

�K�&$��?ݭj�K��3z�����4sXUh��a�����-�k!J-��zQg��k1�p��`Y�ͰM|$at����XH� {g��%r�h{��FX�C����}����h�`�L���IJ���WJ�
M)��7s��̿[Z,���}�-1yg���S}��g�0 /�H�*�R�RȍH��'�ZU�9# ����X��'�b�ym�NA+�P�)���`��?�zh?���{��8�����Lwq��6�O��$n~X���|\[Ӕkn��=4�?$�\� 8iE�шY��ƄtcB��}6����%�����Xi�L�D�0�3�M�D/ϼ�F�-��f����b��.�7�\�

�N���3��&�D� �D����HBq�B/��S����3W�����+�s�}�]L����*B���Y�o���w���:E���Rk����l-B��O8H��H��Jpv�y=�&��S!��"*)��':��2����kW��	2p������c�[��m�yS��r��Iu�GO2�VC�h{K��Pip�p�t�J]ڱ����vr߼
�1{s�@�X�ԡ�����#��)�3d~s�B[9ݎb..�L&�<j�|؉0O�۫:#��Ol;Hx���(���j�_�ڪ�8��U�̃K:N����h�B�~uy0���w�nG��E�U���_����l'��(�X" �ұ ��k{�q���}�U�ᩛ��SSS��<����@i�:���μA��G��<E�ؘ/�sM"�����Tr-�i'L��?�'4��R�3�y�.���a�_y���6���&��JR�h��� gb�\����-:-���V��������r��eZ�#���0oT9��#�����ѵ[X �o�_|F9!a���|����<{��xĖ��䊹�����;@�@�LJ*��.�6Ń�)5b.o�-_�=���W�״�i�x:713e��Sѥ�X�5�s��1~�\R����5���n��E)4^o���;�c�:ZL.���r�ςikk�Ꭹ��i���V�c����trt�ˡ#����lua=�����%�"r�x��\Ѭ����u1����e-9��Cm��(侲e9�ޚ��O���4��<܎��@_�����k�#!;#ؘ�o%�^@�*��]&��KO<��8qi"'UY�zS>�d�u�la�_�����<8���׶v�x
	tM3�+(I�;sѶ�)Ô���P�@���{�]�(gYk����h�	dſ|�O�|g|I��s�����:06_'�_5Dqs�d<G������ʗtB��ۯ�Bt�̄s����.���,��͆'=$��Cj븗��b?�Ln�u�{�|�2��b�m���$���;85ϩ��'���PM��L5��I��?Ύv_K�w�m�]�7������#n}=e��p������6�"�F\���B#�"C���^��!K�SK��Pf�"�%7A��Mt��
�n���1���ƶv�=!Ƹ
��c7�W�X�yq.��M����Ìٯ}��3����i���Ѣ�z�XBؽ��|�?�������lA)��(I����vS(H�e�J�rL�y}>q7�VJ�-��1^�
G�-���V:,����
�iqs���|ԑ5��da9g)_��.#b{��4=��������{�	��6�ȅ�����D���(�3�"������223&�4�@HS�2�����Bv�M]Cչ	��Djs2�Z�s�]�Q9�j�9vFT	�<X�Ŷ�����0���c,S�A��T���72U�Oa^p'Ml:��������*�����Dp��pI�"i6�)e���@��˯���&��8�p4�^]5���xo�F���tp���\?|r���D���V�s}K����z�GP����~Ҝ�(��=��5���Z����<��/��g ���I6��h�s���כ�6ܲ�o�ݯ����qT>���C+�u%Y9���)�Q˛��=5u���E"���[P�_҄;52��F��>�:��!c <��*����hLK�>QE������;��y��W+~�
��O.<c�ݏ�wj�n-��{(����^ݷf��'c�ZBQ�T@���r{%m撥�MՓ��ذ�ھ�#��y.j�C��5�vA�b$���m~$�4K�T�>X@U��N��d��w�}n)��{��/�>���.��*%/$7y�)�{֛��#�D�r|�K���I����5݋�9�.qp� �է@�KzO�>-I�ܠ&�H����S�y�ܰ��!"@7_/�MMO���oPe-�]!0mZ��ir�6"3��X4�#/�AU�v��l�&PF�=}�9�=b��~�ϙ���LM.��ۣG��##�5�Տ�,T�� rh�)X���p�����5s���\�÷F�
;:���Q��2ܬ�열��~,� �v:g����\�>�ᠷ:��V/�O�p��"�yil�X�Y��Di�~�\�j6���&�R�Oyi������m!v�]�*;���0�Kq� P���[n��EV�Sc��b�ge��V�`1�r�	љ^V$K���#��f?�7`p�cI}��[:S(�%���1G!�D��%����j�����綧��Oq�H���1��m��~����Rh��d���p�{��Q�7��7��n�c�o�wdJ��Rmh�w3^�:�:���jF����)����P޶-7��P٣0��#踀���z�$���P��-f����\O�G0�#��JYA����]h���f�S7�Hi|���Y�>\�p�-N�����b�ddأ�d����2�A��:��/��vM^	>�Rj�b��Ge�e��u;m_���;�`�*�@�[<��3%�]Y)4N.����uz�#����ww=�XRKl~��6�q};��k���.��y�[���ΑG�=�7z}�=	�E��;w�CXd�r ]$����W�T���E˺3��}}�Ȇ$��n��Zͫ5Z����t��,�=#��sMaX�>drZ��~E��jp*j��
�Зu~6h�߷�[;�%&!y���QB�-�ɫ'8P����M�ҝe&U��MR[:���
�b�5����*QbO.`I~{�t�bY:�na�ǘ{�]}���J�U{��M�- 1R2����G��_�jA?���X��U��t`Wbh�v�S@��҃է�����nՒ'oH���nv�}w� &���g'r`��x��z�eN��}~�^�\?<Oq� �#���bgM�AAv��6s���I���]�'x�������R��!�(�W�*�"]�	S��8�~K�%��5y�GAMT��s�(f���͎�ܦ):���9�{���~�׮���[�G0s��G[%G[%�����់l��,�iYqW�+�p�#�g�1%��y�`�P$P�d�s�ģ�Wn��4-$��^�	4bE�>\b>�U��/�Mhhg[A:�o��0���hWz[�����*��9w�]���]������VÆ�Rj;Se���(�Lz��?���҉d�/8��(�&�j`�~`΋+����rnG�u���}���~衃i�>`X`��m6<��;���N��h�MmZ~�����Υ�h()O�]y3�rVo�p�C�	b�>I�z.f@=���ԩ���t2ep�*̐7ò�K��h�R+�\��[�ݝ���%��b�Ä�y������=����~�ط�����.!�C|���r\�x���zp�72`6���/~I6rJ�������&�i}����)��:�C�Qs�W��[I+�7�`�_1��A�?رJrn��.�{Zr���<����Hc�D���׻7�cUĝ	ɳ��͍�*0����w�U����rm=o�8���?���~s��,����}�;�W�6�s-�'�.A��!l��m�s�y�ؗ�L�7�l�\I�ѝ,w�kF�`o��mh��Ѷ5,R�x�D�wi���m�Z�=b�#6�v��j ����{k���$e���k��kV������B��ŁNL<��+$���D����1qWK3�V�,�L8�߅(��m�(�/`�IZ�P�ƙ����̒��I����8��v}Ӂ-�*��
8�9�٪�{"����nU�w�2ЍC<4GD�(���J�i��j��<J��o��ٙ5�@��.c4�_���v,x�~�����ۙ��R�����鹺�	�����	�tAH�P<I�u c!Z���D"�LYQhH����I��@+RZ2V��z���J�����蝚�ob�-w�T��8O�y���|��=a���͹��?��d?� �М�<({��F�_`��u���#��(�V��g-%�z������j�y�-�;
2Z�p�M������a^Ͼ���T:�3�����r;_���':�U��"iW�+N�ΉA��lƚƨ	�z� @M��Q����81h���_�ܣ
��y�Ϋ��1�`�>�� %q�Ƙ�����p���d�a˭�K��Ki�7ۣ�&=�5�jƒ�d	��wzS�����	�?Yv����z�E�f���0G�[x�H3���}���q�+��Zq�	U�*C���f<�{S�3�au�&�l&�⇒`/'�@�:���q�A���|�K	�H�D=4J���^PT�Y`��D�O���{}���of�Aj��*ڇb�ڹ<��������Gҝ��U�:��@�>������FLە���V�d����8��GKf6�5���<F5� eBN��;{rW s���4x&~/F�)b*N|���M���p� ?g�o�F���糮�J1ny��ȕ
�K�h4J��n}Hm��:��2���S^ac�!�{q�B��#��,;so�'Q� ���5B����`��/���������6��|#���2�՜
�;o
���|�[��xF���К��A:?�EI�������)�q��ũ���$W�~Ŭ���̐R.�$�:~�p~�\שa-N�[�7���;
�U���w�pU�O�7�H*`��9��Z�a#�v��D�6,u�v�i�f��y����y�[U�yUr����y�_��?�VɆ�Θw�]l4�0#�12|ii���k�l�p�!h�)a�m�^
tB#�Z搪�1��X'M���;ݘ���0����˞P�<X�Q;4G9������ N5�h̽�q�R�;Wr��~wT²����̅��q.�f5����b7��-O�)�x_�iMn�zA}��@�Hr����r�*c�3����f��sH��`�2(w��9�������;��ђa�f��u���F��<y��O�K���)�۴JW;�D�|}c.7�M�rn{�b8��,��x����;qI�?;U�&����l�H��MUu�<�E��Z�X�'<����	��I��Z�Y'�r��KmGA��f��8�|^�N��I�0a�Vޤ������u��3�7�P�'����yX}l?���g��[��X��}�t��b�����V�~"�P�AD�V�^N/�Y�(��;�ABۀ�'N�'*�oP�N:pT�W+	���sK�q*���D���Ò��1	��Z��@����ӡ4>ʔz��/
�^���k����|C��nM��8�7����N��?sZ�5����S77�:)#uw"�*�`wڼ�gb�tF}�b৤�Ů)W�Hf�f������.oy����sH�ٕ���*��DI�bRk�@(i\��^DZ�D#r���(_s�f�8Y�:WY�y���qi��A���/��'�6�s�QM!�3�A�vP�W}�AUN��MF���ت_�pQ%�+����|M��M�7��XVU��[)<"����BK�f�G���Ό�Y��w7��y=�5�=˨�p�P��P�|OuyЁ�m������-EW����&���z��9����9HpAV����a�aDޕG��:.s����TJ�ރ��c���Ԙ����� փG����h ���xKZ�.���s�qO�Ϲ�fN]7�#��R��@�J)�s�����:�qh
��:�������\��\�O5E��S2e9:cZ�������	U#h���3Q���T��A����A]�|������#��ű�bf�n������bI _��41���}V�� �_��>v}�K}�6��;kO8{|gDnp�q���Z!E\U͞3�uU��ϙh��)��@i��% A	q/���t��U]7"�#d.%�6Sn��VL1���0D9(m�$CR��s���?��l�u,N��m�=뺈�I���E����/���W�?��|$~�\f�k~va��Q��E
��(�JT����]�&�n�3�9��(#$1��
i�eH��Ǔ�n�v�9�5l���&W��|]0)���n�N>Zo���[lzZ%�./',>$�.F�׬������ߔ�&����s]��ư��tƀ\5�9�P�DK��i�V���R��\.筎M�kX�EV���&$��~3�B~,N�I�~©/�:c�1�6�h"�I�'vU����g��o����x@��tD�*�1I�a��w��R���UE�W*�I�X>Xn��M��PW�N�i�5�<BH�����ߋ�5�6�Ct�U�b'+	e=��d��eB5�,Ӭ�BڈUR��9�}gˇ��
^��`�d��l?��}�\�1�#���Al�q`�/�N�3���Ģ��6�8y@%�@����m#g��Cc��%�����˷������`Y/JI(�Q�f>6��	��͸Uc�\B�\�~p���|x�+���������D�S�(����k
�E�s~�������ZBCS9�@�K;�`���!�Q�_ID&���$n�4�
ۑ�`Ẃ׉��+6�d�͵%��7M���S���� o$?�EC�<�u���N�v�j<o
�V!�t��O�𑆰���Q�>�y.&71)Ϥ�BU!���=.u-�D��Jo������]� ���ݫe�M�;YI����h�܀�>�lZ�;���X�6c̈���f����yxr��aD$P�z�ʊ��&n���� ��*��Kf������/kA��~��j\�D��^���{���ԌwX�I�\��rF ,�:|��!�1Rٙ����~��Ap���o#�tڲ������߰U?��'����Y^�qI�P���'�2�	`���Ғ>�J*�F��-9�2j�dU��f3=�@t֍9�Ŵ�<�y$�p��jӖ�ܵ\��^g3Y|7B���i_���xJ��h�6����^P���iw�1@�Zs�d���P�͹�G�w��{H�9ʶ����%�M1���_���?�*n�o|� ��,/v�˯��r��\�qU3i5+�5ńo�[*��V�����������-	��)N���#��Ž�n�D��.f��z�<������ϔdIm�a�܄޴O��쫤����o�4qG�Q�J�P&erV��	ei`�&z���M֟9��I��(���f��Hdu�}[�0ź���>4Z%z�l�$bg��gjs@��Y-��ר�g�B	�^o���7.pO�4����@!ta�3�MSj��1�5��j�]�V<2k��:Ǥ��j�?ЌݐK�d.#%���m̃L#:ڕ������[�Iob��{��uP"�[;:~ �%lR��mtq4v^qл�-.a�Tn���d�5e{u�6v��
���|�g�z���\�i����S������ʣ�p���vr�$+wzr��p������r��WM�Y��]~M�-!ǐl���%�?(n�}&#l&���`!D��$�W��S��L��ލ���z���#�,�
<�M{���1�*�p�׏��s���i2<�M�j.�Պ��d�.<����K�̉�nY�Y@�4�BrTת�j�y�1�`ǣ�>�s�D,ICȶ�ф�
���|؆��߈���=Oڏ�]��ZE�K��j%��(~UA:H?94��p��0�We�&�8^�q�֮��� �Q`���%�T�U�$��rt\� ��������ee��]�c��*?˷��*ꎪ�H|
5ܭ�� �oѧ�'u��-�[��N��?p��?6��/��o�~���oG
���6������>׿9�#Pߐ� �Z3��ꥮ-
�Yݟp�@��6��-�/���y���zˏB����%I¹S�Qk��9R1Pp�x('���d{p��N ���=|�[p��l)/ے��K�r�I�{�X�m�H��[��ɼ=�P�M�<�����h����4RQ�\����SE��-'����7�tl �:VCx���s�0�o4���~Q�+.�(�u�h���+��2/����eP�7zʤ���:�y�C�x�ɾ��al�[�^q$>�+�$��ƳԎb�}Wo��^�&�#,yL7�|Q��1��>'�R���&��/d-��e��ݞS���;��ށ��Լ?�K�^p��Up��ņ���AՉFآ�L��7ZU�,�������=WU�&p)ɜ�p�	�V���cH>P2m�>�^{�P��.�}�{%�M��{ji?������tUx�]� ���	��:7��!��jIT=��0,[}��>�W|:L����1�)�˽%� Jx('ח@GI½������Z$���͛ܜJ��<JY�Π/º����@��ӑ� %�����Q�G]a�B��R�C���&��"�咑F�����딮kT_���D(��=��H~FE��� �5�5�lt&K�M��j��]=��M4��$�N<v��^�)����LG4�	��]5K���m��d�~��:�;D���u�W�Qȍ� 1=��xL\'��e�j>F3��|�&�Ξ����xm���(����H�'����*��v[N�X,���7����C��T{������T2ސ���D_D�ꃁ܏��}?|�6�M±��~�X��i�Y]يԂ�=��FN�]���s��R��R}B3��^�'�eJ=��n�����2��_Q[���S8�֓�%_H�{M��o%�2tAa�F�^�rP6c��h��> ��������7f��p�-�Hxc|�/Sb̢f>�|r�����:���x�|!��cK�]R��d�_KD�)K��r���/P���zGߓs�؄��ȇ݊l� �҄���@�çU�V��&e~�*Nk�3��ӝl�(�O�A����~��7>���~k�_���&����	��GX��1��-��Ĩ��R�F���O�I7k���)�ږV)'�evt1�{zi�Q<�{!VX�P�ӥ�J��{������iF���O���!�+���V�6tRh���P�!}Jo�8pr)��=�R��Fה����F=���j��5B�t*��|k~�-��-�\=%I�T�"B��'�s��wG�C������۳�.M]�n"���W� �dC�ħ6��͇}��W��\���+�,�lH�����d�v���|"ؒ���Ʃ��n'��*!������Mc�Kzѩ�"eҜ	!Z�KT�{<R|wWf�J�����@��{P��ygCХ�R�>��#���}�lA��l���p"G�;|���W��Ŋ�Q�[W���v��)�ݯ�L)�5��v��gB��d��]y�t���P(4n�\o�8�I��W�|� �9�������p ثӕ�{(87������d�2���.+�0Kq�)�r�|\]r�M}␘vH��q�[��&�"晐�SFq�>�/U)��@W��f?�H�H����(^l���T.{�S+�8K`���b��pr^�dW�lQ;�::<U�?�^ihH�<�@���0�U���R^�bB��M��v�=*^���'���Y�7������� ӭ�6����'G������_$�s��*�v�vs#+�iHm�����a7�X+��2E��-�P�[�����g�����-��e� ����=K����:c�V��r�͔���i���"�A�,۞n�]�f��X����uhd�{�[�#k�2�zD|�4��_�h"��YD˯��9B9]�(�.r�J�{÷6Mg��+�:Yo���3=��z�N��$��2s�0B'O�9[��������%ȁ����*�覦T�̳�?9~�l&�C�0}%Y�C�_��e��<���qgn�δ�O�W�q[oV�$|�1܎��l�H�pa*1^�.}'�&f9�l�eM���
�R^4ԏ�U�.m�3��˫&a�?��Ix�*<��FX�����d�a�.Ȓ;�\�N*�+},0�JGC `{�u�2
gt�[��	��Z��+�T������[����&��@7A;���<P,P�3�ٞ��U=M2� ;V�B�	EK;���n�V��+�C�J;�Y�0� ���$w��"4��g���R����/-Mb�z*������/}Te|ޒr��pVw`"��H��@�%�Z�W����"�Zuז��aOY�:�9u�J��ih(b3��jo���E�ڽm�J
�o���e���b�d�'U�4t���:�U~D�I#�<��MjG��������A�~#-D:(�L�ԾW��ۿn�k�dy��X�j���;EQ�P��/��U�ē�6vŚ��a�^(����)�
�%��A�zm��q�)}�3bF<r��y�9*�����W�6�M��߆$.�*�k_"��"1�MeH8AcOy�BQ�FF�����|�3�bh?`�-[Ce��� ̎T؜˵��Vy��$X��;���3ᇗ�-6�Yw��2�ѓ*�����>�:��)�^	��bs��)4����<uOG8�������/���v�h2�M5��&��7�N��S)l��4�{m���ԣ���]觖3j�� ��s����/���@C�����2�(��n���BC�_[/�M����Z�J��in*% �+�'
��̪'��q{W��,�J~ji:_4zR۟�Jͽ�m�Z��X�QW��JҖ9��d/�u7��u���hj�P�D�l��Iv!$����T����E]̸��/�����2�#�^m2o�?U�q����Zn��=z.���*dODW���;hZ�&�S�H^8?ޔw�-z�$��I�._-/����	<[��'��<�c�e1 ���ͥ0+���<`��0ܖ�U9���б�Ƌ� ���CA�Ï~`��\�f��P �w�'1������ڙ'���w��|�۷���S�A�Φ��|U�e%a2]������hB�w����0����ҹ�^4�*=!��|v�8�k]V$��3��W�$��w9I�x��D�&L�Cl�T갯%e@R�+�����C���y�n�ԌO�h5�s�扶ӳB5�d%3$��8;��M��;�=�x\�+;QR���-�ܜ/˜_�a��\���d�b���%Yo��Qb�q7�Ia䨰Ƅ/N��t6*y���}%8��S�<M][[��&�<�/�Yr.���t4,��uS�>%d�~x����ji��@��������{���՛t�&�C�Ŝ#j��m��h����;�~����'�^\�ݲ&���o��-2C��2�I�Yg�hn����]D��@T�Mp1>��}��#��OĩW%���e*޹���]m�+���T&v@�^0/���]ﲬ��ut�[hN<H㇉��Сd�>�%�՛��i#�_<+ /����Y����B�n�[������}���sz=\�W:ϓy5�$�%��U8���%��Ť������U���k�(��j�ݿ��E���Z���HU�j`�����:|# =5.x��B��.��Sy����l�z��H`�#��b=��x��"DQ��#�Z��s���������8y���[<4>R>��VF0�<Q ws���M�ο��;��k�~���7M�7��T���kΫ���w<����:2�E䧼�h������p����Hź#9��`�vO��P��+�i����p?b��(�`�Em���n(Ky���\�u��ݬ����a� pD�	�՚��'���K��� �}%��r٩:s��e�9��*��9y٣C`<$����*)`n���6i��c��gc�:���_Ȏ��JP%6����[o̗��z����'Z�<(�P���Up��U-�h,�t2�[�~��!�7�Oq��M
���#�@��N�k@}��9�X���
���k�y8�AJ�ʙ՟��óю8���\�}���L]>a{l��^��n����d����Fz`/��ma9��4�?6��A�X�f�B�y�B)��WU,�E����P��6q��|�~_�f�����m�Z��A�Py$�����8˯,*}� :��Yk=J��ҍ��g�����56?׮+�P�����	�~�AȄ��@$]`	���P������-����{"��?�G�i�����Y��ʉ��>JxW[�c�#z�+R�]Ft��\�ͯj��|ZU+ːoO��'*b��}�3������5d�����+���^
�d6cTܪ�8ּ
(,`�		럯� F@Ԫ�,H��hmE���ߺ)#��a+�ǭ�\KZ急�l�����ߏ<��l�M��tՋv��ti�d�(J5��g����t��oy�2��[���^Nh�n��w�>��{�i��+�rDժj��q���j�7t��7�b��-�c�ڧ~
dWV[�_/���sa�����y�ގ� )Q{��*k��q�H�n]s��-R���-��D�x_4�����%��o�t�NS�������`o���;��U �>z,I�J*?�Y�G�W�i�zኺk����Xp�*_C�����b�����	���*��K7"7��f{F��^bI��UI� ��\��S�׍A!�ԉ�!� #GD`�5}�w�L׬ڣ�sy3��� =��o���a���,Io��[� �҉�_A�������T�#�'���z����Aav����SVlM�z��� ^yϿ5��D�V��D�I}?��K����oDu�=ءd����r$�\� 59�(߶T*J��fO��W.�
J��.t҅���У$�1��_����<n��~EC�4��FQ�W=�pzz��j̺>��nK�U!��%��Y�Ω��8�%���˚;l�\�T�>U��H
uÇ���#���É�^?~�y[Ki�WA��Pw�i����f�t C����lF�x�ߞ���h�O�՝���Uo��u�V(Rܡ���C���ŭXq�]�;w�����z��ߝ�g2������k��J�׈r�|{�"��쏞��o��/S�Ѿ�䛊��X���U����A�Po��Y���5H��2%V��3z�B$�l)�����I��;����k��j5�iS�Ǵ�.�ji�j9��▰W�o�:Yk�W:֥n�:X��H;�B�ۈEz���E��&�k5}ҕ"�H<#;��(a�����ޖ�&�D8�6G��9;|_�f�k�_��kS7@$�T k�Hv���t�`�8��w�]�:7쮁a�[����J����\m��r'O�w.�k�Ȩ�P�xՅ�ޫ�����Cwl�~�� m$x�����BHf�e�����:րi��qO����Oz����њq喾�=}���R���5r��#�8�^��e֪��S�Y`�1=��	yeeZZ�9ƹqM�4u��[0�K|�����(��[�<]�(���I�M�G���ѿS�����^�【�g����Ɗ3�Q���]��ߦ7�7��g��l�D-�-��1� t.Z',��2��Պf���/a��ǰ���N9�"4P-��3j�l�v��﷗�j�5�:дE@�Q�?4P_Rx<�>v�����BƸ��L�c�)=x4�$��H�[#����
�g�l���)� �/��{x�Ң;�-Io��q���ז{��v��f�g���1�[��	,�b�@�y����p�E�GR�uV��z|v�ldg�����w�6��P�u��Ϲ�����Zk����ǐ5i��q�=j�^/p��	i>_
���a'�ka��߮aM�?��>�+��d��R��`鮪��6g�;������Xp���|HCwU����c��Lq�ٯ�O�ܛ�6����Չ�T�Ld�YMn��Wޘ�q��r����_��%���<���"hwp��Q�(��BO�_̌}��makh���QTU�c��*T�<������&����LS�KmP<C���=..G���ݮI��L��acC��a�L��f�e�H��XoO[����Ewi����a��~�y �R^��.��b3^��u��@=���_��߆�@��3G�x�)C�d�;<�67�`�����ef[I��6_�X�8��?̖��/���v���.���i�FV�1�0���H�p#D���'xP$�e~s� Yش^���ϻ��_�:����]�1���D�+dx��]����rU3����A%}`��F�u�ju]2P�1�V�ߩX�4�@����������ҝtg�c�,+��N��A�JQ�Z�*�["���u���JUe�;�-#e��-����O����ڭ[H�I81 �,>}nEX#	D�����g��ae���o��Cr*�i�U�~`:���Ӑ1K��hRn�Ms���/�/v�8��,V_t۾"�f���Q�C5Eee�'K�q�h~��7aR�}[�E��#(SUA����5��;����I��UQ�qX1����y�I9�1����[���-~�{�!���7{G�`�1r�^��eD��Ɨf���e�}�J���ʍ�~ͬ�Y�G�o�:-���Ս��6u�lB����3��\1�*sЕ[�-*�����[����_w9��q�{V��^]�xrgC���?p/I�4�Y�����'�,Ci\S�>�%�~���+8q���F���#��#}��so��NH��9O[pD�ƭb㔛��El�(Q�ߜ��f_�)ů-̃3�UȪ916�k�\w@55�/ŪX%�/�L�a�tU.gzx��R7�dɞ',xzl�m_�I��s;���b���U|�[d[�'�6������*8i�:��%�~?�)0l��c�Kog�E5�3i���":�ٴ�d�"�m�ڄ�<ԍc���I�ros��j(6��$���z�����1wl�~��a�j��%l� j�y�m>؏�*2�'�[��~&i��h��y�@��Sӝ~�h���>�W�<�����M[(0�g5�=���6���BX��(ٷ���	�^�o�����I��6I��B϶���T�������vg���,+�,f�����U��y�`Iu��5���c	9�	�nݴ���(��q��M���x�ϙ�u����>`B� ����mUa���_-_xr&��)��eD�S��[&>
����|[��^0Ll�Kh��u�!��k���f玜���(3�q'o!F��Ʒ�'�c��_�t�UK)̙����C����|�»W(�B��u3��V >�	�8d�{	.�U�,Tj���y~��g4�~DJ��'�aȵd�E�N`*v]&ᔙ9�,��U͔g���2'��8�|C�gR׶������ LY2��v��X�N@@Pm9G�y9D�nL�+	S+�T{0.�E�~ ����2ôy=����D^'V`����.C)р���Yy�ƴ��H�T�H��-:=�nɌ�n]a/�X$B'~K��d��@N�cϪP�_���z����#�߁C,�XϷ����zneIFb�1����7�����}#��I ��i�'�*��U��!a���u��f������ij��mhZ���7��yI��dx�&."t$�H�H�� Բ�9�m�7�,�k�TL
]!��)�F:R
Y�2�9�B�/�����+�u���Aqyy_$�:t�#��_�+���ő��r�LUm������L�	��p����Svpȟ=�SH!b�GD*�[�|#���ض/����\Xx淳Cw�ϿYƃ��u߳�����W\tp�))�5�>���;m�-�W��6�zC���y�_����0����N�Vs�>c����AFH�!��9��Cy�x�������ۢ�WT׋��@�Z���h�vaF�W�?Zo�ݮ~�Yj��.��8���"7]c_�k��V�=!�>!�o@<j�9�آ�1F#���c�x�����8�f�8�ư7�GQ�G����� ��Tr��q����x/F�8t��Vy���*��k�;Nz����w�p��\bfcM�Sko�U��n�V7����J�jVv�pt�?�)ָD���n�\�o\/-���:+j�N-��J5��w)�:��L�W�-���I�,:��k�e�Qi��c�6�K`
�΅�b/g����UA���Qwy����C�d�^i��~-L�t�nX�H�T>��3~p�.�_b�mŸ@"d��п�Nwx$���5�����ǃQIP�������=�of{f���@a��RR���b��c#�\� � Qj�X�	Lt��o�LI��!�N�ZTy�]�s#�'zpQ��'����Ᏹ�[v������[�ܟ����?T��l5Z���'|��Ϯ��ȴGH<�߫W�E&&�L��ftv�i��*�F`:QC?�X��i�Iۯ���J� [jZ��y����VUw��� l�r���8�c��͆6�<�8"tы������̋�:���ҒB��쾔��1��쯟�|#~_�O�����8zGB��~u ���,��N�<oH��fk�|j�3��a{��ß|xu2�� �U��.���[�
���J�8�~�|�C?c����z],&:��_���?Egyi�շ�HS�c�QclW��y���4��Ђ�O�s�Ǐ�_�ҫ � ����`��	]�#�+�*�h��Oc�V-������ m1���5��ZӦ�<,��m`��r}t4�/<.�W��õBN���T��T�����d���:���F�蟧�'OHl1*QH����\h�Oa��U�����Bv&6���Q���q���(�2���@}���Ϩ��w�ͫ���x�끫��:��8Z��������Iw�/A鍺���,��X�L-�!J7A�t��p����1�1���E!ť��,�a�M����h�� aJcJB�Ll:u���5���Z���@̖�9�A�Z��Vq6>\�ff�v8St%]A��}X�k��78$�2�Q`*H� �n#&X�̹����O:��&���,��Qeyb(��ě��N�ھy'w��Fd�J�HOYy���_]���`O__�7�7���?�ؔcV��~'���6]$Wգ/+1#���Y���N�YII6�bΎT��������caa�����T�j�|VU���{��>��e��5�ڧ��}6�##uV 41{�0abW��������� �rE�()ޱ���1��{�����T�������v둈����@���rE�#�m��Λ�pm�qsjb�p����̡�`gb@P�DA� ���*k��E���vo�	=���Z_������"4m����Y�:&��i��|�m�%}�*�a�$�;��_1��ly����)���5Asȣ���臒�(	��e=��D��'@{@���N��m�A�O�]g2��[�T�m�`'�Ev^۶o�D�M��l<��Mf�ps+\��T�u��ؖ팊�rlD�^�;�"H�:�#ۈI�3F��)���rJ@�O+Z{D�������O;|��y������/zM(��֯�0��$(V�7}��h�ЫW̦���D���>���̪��Z7qW���H�Z�(ԁ�MN���㡡�X3K70�݇��������
�t͇���r-Dy�'FH�1��Șa;�[F
��ó�{5�xM/�"��:��a�tv��r�]�-
�#�q-#|��
��F�Β�\���*j7�=r�G�$!E��C�i��Lp�Ӡ�	h�[s�+ ���֢Lh�8Q��A���(G���Ä�G��R��,$;����3v|V{#_Y0�t;�-ꟃj�=��V������Տ�>��(��$1����!M��2r���i��MC>���\�Ș�<}R�-)�˶�P_�Z��	&�^,n���>��H7�I�p����:�j�Ս��������%�;�H
�̱GCJ�\M����1�����YQr!�߽MyY|�{��)�0���� ������C̱-'�JH��B�"׷e�v�FPL����(}�:%A�R"�_n���5T7���	�{�J�VH`��ǎ�`�.YNg�Hlo�j�)�b��5��w����@�w���S( ��kA�Ί�Ts����x��8�P��v찵l�� ����gO�I_ǈg�:(�Y �[���������`lO��<.3��76��9D�5���Y�����V=���_�|��n+v�.���Ș�~)U����g�5o�J}�"%ƻ�z%#��?Q�D�6���8 �U߇l���(��_H_�sW4��vfr �bE����2��Y�0:�=j|�R:�'sPs������nL����"�G6%�_U���@	!��3�M.-�;|?�����.�w+?I��N�*|�j:�q�0�2}W6�>�x��@vGvf~Rh��Q�����,1��`!b,[ws�R�W���w_vW4�r8��'���|��HUZ?�q��G8���������C|$"Bh�g�˓�Ƨ�eN_.�<�Ľ�%�#�t�^���]�c!fh�B��-d�~g�|�m�!� F����jϖ�"���~���Q
��[F��l��}����;��ng�ʐ��x!�6��s��(���@@�{dz�F�D�Xp8�CU�F��kd4_����9����U�ݓ���U٬�>���ɏf���k��o���%`����/�!���G�b�p�m�+#���{����!�8I��-ɤ�=�&sL2$5&*;��2�rdf9@��s
��Lo"P~W�J99�Q%�x:�s�O^��_ڳ���9|9��D����_��<�6�9D�u}�����*��	��vMpH�ϵ��J�b��m���7H��9�
���|��;eF�.��=c-�z�=�~\��a�E=��5�6p�,�ujz��X9dEl@�	֪mE�bj(ƶn��d��T��Lw?���	�j��/�A��@�[s������8|��?�K=�0��!+P�c�#�?Q���7�}�G��e|&_�\.k�ި'�Q41�tnmi�%�X�׺ :>�~g:ml�/;C��mD1M�`��O7��l����
f�^(q�2�~=��8�-3�;��d}V\П����t��Y)~ƿ;�4��~Mm����d��Ζ ������($2�w��{s��XMt���\������$pV�d��?d��0�n�+��������h~��dw�L�\j���2��6k�����J^Ȣ�g���Am����9���ȁ0C ��5�AYmA��Ω��ʎ����6�\3�� ��b���%�.���\�mG�R��)ύ ����S���j��zY�����jY�:����Wh�K�j��H�fw�í�>�3��.�¢�ĩ ��lJ�F��P(�h�cP��`R���"��(Ivh]�N�vs�D�9�6�8׽�t��e��(1�M��
-`2��*�kNSh;���(�#E��nm��`1�p�ЏͫW(�`Hv�6��:? �HT[� ��e��b��)��i[���4q��-6B��)�˖�j�+PZ^�����2C�-���̘���=�>���Ft�����k�6�`d��sb׬�Aa/�Z�2�K����oKO�\�al��f���	���2�9�8�bЄ��v�1����I�� �W^ߥL2~Mۋ��}�GgI���bI♖��-3�n����n�gffd�[[r�gH-�>.o��uR㻙Xm̆n�籓+��V�:�I\��^�Իo-S����>I}�� �N�z�|����?�QZ���ME�]Z�o>�8�T�AF8R�d_ɜ]X����Ĕ�(~#B�P�5�l�`���\B$�sx��M@���_�ְ�w�S��Yg0U!����*������3���w8	��66�a�~�y�"AH���O�kPz��#u�a��3:{��/�=��}���hQ�u�P����yQ� O�;��p�n���n�L�'oi#{�o�ĭ��`�m'���MD�
纟P �{��MKӞA��6܌�0�_�d����4�~'E��j�����?��:�%C͊��ј�1��߶�*:���N��ɀ��nͣm뙨���9�I�	��8��$8��}^��u����@��,F���M��HĬ�`Ez�D�s���W|;E���+3(�bN@ �%N/tB��L�W֍��U��}����ַP�w��0��$�c�GW��n"(��AĬ��㸰>M:��Y"'��>���Fn�"��e��>�X�?�P̓�����J�V�����Y�\A�'�˝���N��/�1
:���\Є�~�����B��sZ퇿��<_�e�i	
�WT�{I�9�>��,�l��p��yB�>6����{)L��T��$�2��q�ֱ�;'�l�;��u3��e��5<�øl?�[_���
��v!�h��ѡ�^RU��a.fT�r��L��w>/�q`��DL8v�Kx��/
���� ��|����r�߄�)΢[��4p�ɥ�{|���%)��?j��~�]��K�^ƕP;�r�5t��3[WT� ���-���b���łd�ρV`k���K�L\ǿ9� Uk�Jɘ�"����w�_�r��Z���_��"���}�����A�w_@A�n�c/^5J��5��(�(����������Cu�w8"wx=�-��ۜ�ؑ��T;B��_8��a��&�Y؈�6c��UGM�/|��M�\��<��a"ɒ TcÝ݆As���l$��]_:���)�R.&$e7�V��O�-I#�������?�9OΫy��BV_g���$O;
�k��|Ujr�)"�OY����T� �3>�v_��Jky�^w�ܯ�d���t244|��Jv(7����X�/n��ao���%�
�/=�U`�&a� ��EN���Z3�L�����V�f�I�RM_�{����ĕ2��\�g{%In<K�[�T����u�w��ԍj�ܫ��f�k�b̯��s�'d�]ɔ~��zb����9� �JI!1�5{d�Ϋ;��L�Xq6779������g<e��8�8�-��|��UX��٬�i7��w��n��j�}|�~�\��MD�n����K2�>�2��^h�/��o���U���:�� �a���ѿM����	�-{���Q�;��Sm��	�,�2570��5�t4�Z����e�$��Y%��(~Ta�U��l�Y�t-�+$���&�8����:h!���^����R��^�֝��ļ����[2�[��z-x�ˎ���3����
��ZΌ.���I�lT(���?�-�a4{� "�_:�C�Hrn����:�����cƎLgv�~�21G��(�"�Mt�ԋ�TI�ʑkK������໎R)Pga�9�?K���n1��Qb�Q����p̯e/W�r�oq�Mrd0b�:P4�6�6Y�y;mdd��u����@�⋮;�M�׋���Y�EI ����wz�� ��̂��b��759���%���+�%0E���y+;�Lb�_�h�:�'n�YԐ3����8��l�ػ��i����,M�Y��ʼu	U�[����޴ �z��˱�qw �O��$˘%1��U�=Z���KyIs\���a�AT���q�K�U����O�����4E�@�GԆ�W7Y�Z�v�~�E��ь(�t ���\-v�h������?��oOX�� 2}d$+��	&^��S�
z���W%��TI6�ݹ�Ʈ��B��]4{��ۚ�������M_�u38��Q����^�X�NJ��_ĝǪrCm�����Xꠧ}'���
�����MnN����5�@�к�S.�1�`H��*B�����q�V��PR�p��NY�"Y�����%���p�"pG�ر�"����,o�$��|vz�?/��b�����S���-Be�4�}��C�l0�^\�O�˝�|(~:�<{�8�w��E�SQWJ��i��e����#�F����e�vg8S{H�L���垹�y�o[��גn���>X��_e�m�ǉ�E��+�e8�,�w�e���D����9�N�%���M�
�Xg��tG\&�����:���S���ZwJ��`V5������`���(O	|�SV>�n�Fuj����l�t+���gt���;#O���6���I)�Q��*=L��7Yt�L���������E���y%��?�;o�9!�N����ּMvL^�S����pӪ��7&XMD�G�0��#����7�J$����}5�^O+�V��R&�b���m,��\+�����(gV�<ɗ�q�O�h~[�?2���z�/t1�)��AeX�U=��q"7v�b�L��ܱk����}6ӷ�Ӧ�dP�s�C���J�%�xv�_��i_R��Պ�x� 4��������9O�rz�?YLa��F������힧[1=(wӇ̹�[��q�Xn�_���)���gq�E��,<�����zP[x�_���(~��#u�����K���?,��������o���鵓��rp;���di�6�uߖ�,��i��'z�_G!J�&Z�&� yO�c �-��C����O�����z���@�jd`0��f�'���&ЕK��L� �M!-�
Ǻ8x��б�lW�ۦ|���$}����`8>�Vv[/������o�a�)�j��ʐk�p��ݷ���UYYu٬�mi�s�!�i
I����NŒ3m�fn8����Lj�r���?�0��=�����0G�����v`&΅�.�~���g�"�n��M�`����WY�.\�I�ę�p�� e��v���վ�/iLQ_M����d�������b��%��U��oD���(�e�1�����oL���9��f�\�FV�`�pJa8�[�R��-��������!|"K]��*''��݈�R�a��STQiN|������p.���]q5�|�¶bv�Gn}�t��������z�f^����ǰ3�.K�H�g-���M
�'*e�*I�̃�����X����Ј*�(1�7~̲�*�0��;}H4fe�z��+۞`u�������z��2�d�b���}��b�;�Y�Ԑ��������vr6��%Ec�j�ülb�vGC����Ǫ�~G����ᇫ��m�i4�H�����&D�)w���e
�!"�H�Kϲ��%p�8��A��Wv�C	GC�w;�b��r'�h���h;�DزÎb)��Oϼ���:��K��<�������;m:�,A_�I�9���J"���}!�I�i��\c�a��G�eM`׹\��F�J<�4�c�O<����`B)g���.m�T)��� U��L����R(����a=���H��"��`�}`t�`a`�)<�F�}A��b��Q�dU�̳v�e��;urXڢ��9�ja�[���i냀�f�ՊLK �T�.EH��0�_��mg��M��Os����G`[�щ�%���@�A2�y�����M	zD�Ik?3$��vK�X�+ևx�J�o�,4�M�Al�y˙>�᧛M�t��T<E�C��tV�yl�gx�/4��(�� Dc�`"o������x�]�$n��Y�'\��ci�w).�,Q������m�4����H���UZ�1�gZS�'�L\�w��H:</���� �=�_h�R��ZJ�$���e�tM�y�b���{�"���k�M�@�_�t��,�S��oרC0��J;��H*��6���A�UW�<>��Xl��U��t�_ʐ������/�&��U��x4�Jo���L�OҀLl�E8u�	]y��v��"����O��Ih!h���R������!=ɫ���.T�����=K�
����E�!p�>��aY
��V͡����1�P����4?��� i�UB�lZ��8l<Y��Qt?!�^�<1���	}/b��r���M2�m*�k���F�X����-0j+d1"�ܴ���F"�k�;,�b��'�dZ��f�V��0T�Q�MD��JA#�#�&������m�wg�ղ7�8G�z������n��� &-Pd�^$+�c���q�W����1z���ҭ�Q/��.�?�`� B�G-��:���D7�*Y���1��RJ��V����ooS���?��$���o@�F���;����˽����������"�G6�w�p��Vվ�Z���HT��¯Y��iY0�%PBŁ��J��E�Fh�Y�T��D�����9��ߺ�n�z-�J��P��`�5��*I�i�<����A ���������eN=�%I��'��n�vi��Oլ�7�/M"l,��˶�5U��cʌi �ϗ�������K��ԇnQ�oB�LD�Cc(�%���i�'��L�A
���a=A�^A�z%W	�{\b����-��)�F��튫�y�y�ؤ�3�W
_�ϐ�˧e��3����K~}{�̗��F�6�Dr)z]�ێ���>�@`�V����I��E�
����[�/��Q��Nhq>s���c@L���[��e�WM��&�K5�,��5�8:f����L�Ze��D1H�Đ�VS��.oYh���m7a"츭;����-��2ޓ�Q ���hׯEgT�O4=�){C<���a	8/�$XTm������R��{��oU*=�w�~��-|��E�p/�1�%dE�~j�}�"X����@L���Z֒��$�)�����w�hT^��.a��:޾+�|3�\}E��J{zߕbnYe�����%����u�d�zY���n7>�a��M��u9،bs��������qe_�ؗ�6ܝ{�bc�X��y���,Q��5����~�*{j��+.�y:P�R�~�����4%�Xc*c���[�?�Fݛd��g�!]"���*
�y^�yDab��?&2ꆁ@ ~���6Y��%SŔ���Zj�j먗:��^k�LX���ΌFd&��(���"ȑ�&4�N�V//wn�X�6��"����p�2җ泽t2�F��D�-�N�R`y�h��C���&��B��J��\�p�a
Г�qJ']"�@Q?#Fܞ�y!ń9�#�ȣ�ܯr�g�`"���2b�6e�N�}eK��sU��*�HC�{\[`JN~�S�[����wR�2�e�I7�&���N�ֻr4�9�|~5��pꕼ���Ld��e����e=�X>ۤ�e�D�~�ڒש�3�>u�Y�iA�x���Ț��Pņ!�f������>��+�-�<-���~�C!�3ud�zLM-E�&��&m,a&�?~���ǭ2�K���sjx�P�Ƭ4�7l_�5#ܽ��}����`�xI@�7$1N=21w'���ik8�a?:��o��)t-s�M��D�F�x��Y�9U�ґ�c�G��*�]n���f����N=܀=�ݡׯut;B��*�:|4a�r�Jv���m�z��d���}M�)A|V��%�ޏ�.dD��(�$G{��C�0�����@c�ckfCm���j�,�q�ؕ��ODW������{�xyʱ��r�t�mVC�Y[[�>�["�����e�rDI�Lx>h�f)b$�
�䄸��P�P	H�Д춵-��JC�@���H��~C�Q�K�2��Y�N�� $�����t$NC�b��i������\����s���N����!4��\����]��K�b��C���;jK�9��e�0aYz٫�/b\
2�D����ܦ�V�	T5J{�d�����"�L{J� E��&�(��m
�I��H��ؑ��_K��5_,s7/���M�*i���-M��n��p�(�F��0f�sM��^���W`	���ܵ(��!f���\̜y}��Y���������.�M���H�y��Z��r���P�3^������×�c���|�U!$��DԄ�]C�����k�Q�T ![��܃H06����5m�v�?��?��4:��{ro''CĨ���_
� !�@�!h���D�*�b=��}���:���v�?��Aod����1�*���p�t�W��6��W�B}���]�Ug�#�@�X$�n{�B����'�����k��Q��L>hkJ��Ǜ]��eљ�.���?�ޗ�ds�:���,�V��|�cǻ@�0ٖjT��&�L��ɆQ5[������ F	8�:޲��~�"Ĳ�HEnFu7��%&�I� L�@�(M:��S����W#��A�h�W�b���M�$D��sM�["[i6f{�I�ZkLo���H}��`^�Ĳ<�#�M�h�b:Ҷ�WH+c湕@�L�Dn�K�m�٥�����|(����	=A�Ġؿ��_�k���DX��`�p��9��[S1�7�Ǳ�:֛�^�.�|Tu��센v	d���~��� �|�+�_|h0ڹM\t�!��Fex"����5HO�(�~;1`��M¢�A8��L\�y�����>)���yg�3Te�Cu���nЅ����ں{n���#�Թ��q��Î��h�=�>Ky�X&�h�W����cIb�ƻ�J� ��"���`8��m�(i.0A(�@j��������vͺ/�+8�0�$���a�M���3Qڪ��a��t�/1�i];W�iVy�jS�&����E1��*�NU�2����.�����|�E��,%$�6����X�^�G@L��sU����ep>�T��+ڊ��/�O����!f�J�Q�g��c�W�UVp��s�N�ׁ�|�(}��`q�����C,^�د�<ܫy��?�t}��7W㟲~^֢���{������>�8����DLR�*�ΟTs|���,{�w�Ͷ�TZ��]��@���q���F�!��h��^/��߽��k�c�$����[GfNS%��,��_���b�Zj�т�4�$�Q�����j��>��?��}͈�lDk��)����|~���0�uob:���.�������[���K��� l:���v=��mۃlN��2Z�k�>����d�v:��c��GU�t��j��]c��	�-7B�M7����?C���pl"�yK��QkM��jO�F�G� �'1b�=�I�8A(a	��O��to����yxZ��5n�o�h�����d��)P��+���|mu?<�Q]XJ��#��b��$�V!U%1k��	�ݻ��lL�`�3?�,ME=>>B����;�#��.����U?qG���c��/��������������Z.kr�*!��$WE�X�[��ۉ���qm�oa��n��[���']�I�AYϻTй��WR_�*	Whuw[�#`;�`:��Ѹ�'p��Lu�9����;&�
�x���F݈�����J����$9��]�$����Z�A^n�il�0~��0s�G5�i�ʻ�y�ϯw�k8�F &��[��n<��M9�s���cQ��(\��0-ڣ.o�9q��(7mh��,0,�!�KաM%�0�-���$���j�Xv�܋S֪��w�z]VQw�9�ʧ�U�p��O�U<]٘WR�w�4ef�'���4Zpo���J�?,c�]�gX��{��>��}#��T��7���
�LV B��%0V��?�j3!>�D���a�k_c�eHs?v�g�O�&��7�$z)�B;��T�������~����I��k��J�Iݎn ��xa���c`F������m+�A��|%\v�d��5F+R���w<���t�"���\�{>@]Җ�!p�\ť�
#oC@��f���3p��B��L�L��d��i'�l�J����ٝ�d�X��G��H��$PMr�69��,1`���Q  ��������oO��9�p��8z$�^l�:�}*K*��{�߷��?��6��ǿ2��:�~56�D�8t��[�N�b���a�2�9@��
��H�@4V�T���7����^�W$�̢t�&�����_�
1\���1��3�xt�Q?�D�W���r���p&(FO..&��9�z)�!>��0F�}uɺ?�?�o*E_�{���1;ܫq��cG,��,���R��`�XII9���a[���-泤eL�K$)$Yl�v�&�PR���*7G��W��F%`{��whr6T��q�0��T������e�+/�~M�D�Ғ�ko�eTb(�RM�ț䟿N��F�]2WK�d��]��3`l_{E�r	y�C�;L�p�����m��FT� -!�7�"�n�_��ַ�h�E^ΨX/|������2��������Q"豞��%:
�)��S�Q9����<�~�*Z���M�	6�=��_B�����͝�ۉ�4�/�Ҭ3WR������7�@��VE��?@��ܖKq��5Y�t�:�<	��h�F�0���&��?��XG���GT~��w���Y����w�?�~z��l�_M����ۏ{�O��^lbVBt_�;a����/�B]~�HG�>�	w7`"���ϭ:��[���j׭�+���׫���紋����3�4�������<���*�,`��_j�z�6m�u�,�q����
x���P�+m��r���<���*M`:���f��D���e!]/>h\���I��/vO��Y�������BvK)؎��Y�΂�C��M�]jgf^����W+:fM.Ic����p�a�_�[��8�}��  ��j#����7� I�[�*I����L"⣣#�#fU&��^dMB���L�*>�L��L��ZX)��N��|hjĎ����E�4?�C��.TO���ȘCm�-F�0Ϋ�)��]�C�6y<g>ĠPϷ�{l�MW��㠶2��w�$�Ƥ_�+�88��V4�V#Z�2��TʢT��U꒤6��a��7�8�� ���ˉ_5�$�!:=Zv�_w�T]KΉ���_	Ձ�hj�k	X��K.z�T<���;Ey��Ϭ�귍/o�ȡV��0���^���\V�f�krg�b��t���aR�����D��ڡf�.z����@���j*d�Y�h�@1QnBvs���HO�����s�+F~�Јj`����8�L?����@Щ +����#��+�dP�x���i��B[��IB��8�{���纞"�/G�ɵo��K>�1�i���P8�N����eͷ|�T���'�Ef�f�֎��|�7A ��7�����t�$���x�"U�:�#�������~��μ����&���}Q��g��;��*���$�VVP�aݝ��xz��<w>��ﶌ��Y���,����b�jCz���+���+B�q�tNU� ��z����]Ǧ�6��`F��d;��������xٗs���}�*i��W󥹸N���Fd2�f�D�F�B(��O{w/���{�!�vb��k �[�zW8�7��?b���u=,?�D=�8�V�K��l�K��}�] 9P�PIZ�8{h�y%F����^�UcZ��E�����瀚���i<�|܋3k�h��C͙>8Ѓ���PZh>�B:iu{�g�% ӈ�#�I�4�_}�����3���8��ҵ��ǫ(��E>a7Kd��N��i>��cX�r���}X�(Os�\��{���lH�zA�	;Z��L�šE_＝�Ma�;����n�ʦvx��o�űD�
w�i�Ǟ`ԁ�vw����}�JЁ�P�ջ�S�$����:��S��̪�����[ ����5���{qkq)�Pܡ�kJpww)Z�%-��ݝ�,����{�o�f�@&���=g�yvՇ��ً�ӡ�A>:.��\i-ч�������6�~�>�|#��B�u�{���e��u��~a[�������X�Kpmwi�P@�<�_=5]����T���%�Z%�h'a��+Sk{,�t�>��z21�q��5]D���B�/&v����g�D�|U7\R,�S������|���';��
�R"�{8 �z��4���z�~j��B�^�-ϊ�f����r�g+� :�NL鱸�G��h�q)ܳ���k,��m�C󂧺������mҏ�P�`Ņ�m @-�q�T;@k��P��B����u�O� ��/�#���%@ɻ:ߖ]+Y�b @��£�
Tc��Ƹ%́�q�r7�h?����e�:�dP�7ֵ�u���{��Ġ����:��OҤO�$}d���-GF��]�u���R@�W�����wZ��PB�3F�m�?$&��^�"=��* ��?��!�ġ� /�,T����:���&���:Ǜ���]� {Lç���@_�a���P[&�쨳IQ!iȸ��?=!��ݪ�eJ�n4����?J 'YY����_<Yxb�bvSu3��MW!�:�]�W��X�[VP�E=\��f\.(n�o�+iMdy��F����X(�a+ÑU_x˔oR�f2�EAj�%�<UH�Ǔ_!o��$;�����Zi~0����'� p��%0�X�'-2jo�_�&M~4�#ʢK�o���L҇#y׻�Kx1u-Ͻ��I��1�^n��mt���6�solQ^!���WS_+n$���T���|%6�)'�f�:b.!�q�2�ٰ/;>;��Z3S�~��3a���M�b�����xLV���#%���ZD\O6mmm�+;=�N͞�*�L�e��K�oc�a�Q&�]���n�����N�L#|����p��beh���)�7I봅��g�;^��QB�K�a=N��}�}c��n����!5[�>YMw$�@T)�~M��Ǔ��t{W%��&5<o\V�;?Op��˱lFC_^V����bk���)�o�Yi��������a�ҭ[���6�y]��VL@d~��4'�h��\���4 ˮ������f��k��*� (rI���ș�H[?4�%�k�.b�q��9@�,�$$Db�Ͷ����S���c���?���x�F�B�4hs��[��b��c��fA<lZe�]D�s� N%*����\��a���3��-2�O&x����F�bj��XbA�{�ի������G�c�}�O��(�J�F*��=�������^�q��毋����:j4�m�߼�/=����w�/1�w�
��7�J�`[��b�8݊���\v<pW1G�\�E��o�`�v�eA_����L[�h�8{�W�p��?�pt���d���@�3�'@a
�5���<��	1d6.F�&ԨMYt|��ס�5y��6��<�Kͣ������+mF��&$֖s�~�?Tl�u�͘ޅ�U��dj�ߨQ��v�T�{վ��;�`J[�;!3"nB@� ����E��f��U��G�AA!�j/�Ȍ�f�5-�g�n�"}Cң��7-�R�/?(��/UfgcUt��,V��}���?h��~y�����&�
�qC�2�4�9�~t&5.߹1�q�%ϨLY]�����$��p!�wc��Ǉ��+���U#pA���Ô{�2g�0(?U=����ވ��4x�[�t��<�s����v�,حLH�s<��vv���;�GM1�晭��	���#�0H_�Lj�ޖ}T��`S[�	�\���~�6���_8������R��	Q��f�Z��Q�/d��1����7�}�-�\/K���$
x�T�=���i��ϧ;�Y�y�e��򰆽f�W
M�q��;�_V?�'���q|S�F=9����X򾇺ެ�Pzi]����:)��~�_3�#�q�fX�5����� �U�k�����*�N͂�d�H�#����H���K��&�I�����+��W9N�W�
��ڻ$m��6
T�����t_�K�V;m˔��3OV�?�#�y��-	җ�c�-q>���8%[�5����հ5�񦕷���Ŧ�@���[�?0�呴T	���)�d[�E����NE��Yz9�_k(���m�^�*�@$�҃����s*K�ʁ��³M+K�Ll�R8�3�W�~��}�X�G��k|C��mAq��5���@)4�[L��U&�z��#F��aJ=ת�L��병O	:�[�8]�m��Ǹ��f;����ϪY�nN����ݵ������-)�H���������-;,2�\�w1�YJGG'7B�,g�[�_�{�D��YT�#���<飂��H�Wu�N������z�`kRO^(�`g�#��6� ��\o�]�ջ-
�k(Ǹ��=�-1H���\G~��*����+C�{�W3m
��#�\N��C��t�[�U�1<)$3�f����\��y%Ve�絫�N�H���OW�J�6��izf�x��V;o�/� ����|nl�7_+^׬��n����)�ՃW��8򥏂�ҍiE0��`#	�غ�^k��a7���	{��=n"�����nK/m0����k�^�!q��[7�)J�& /F����TF�ղ��p#n1_�Ga���h�2̃]�b�\)ac�m�Śh�Z����H�@���G�beת:��Շ�@U�)X�x�YUF*����Eh��B밶=���=�(�N�E�������L-!Td
c�5V͞Yg�3��@�|Ar����o�7����uy�����R(��^$1��K����~����˥�:R��EUv�ǉ!3Z�����9}��7�>�Z�FR��s��s�C)#���~�m闆{]Eq;�A1���z�;n�Q���b2���A�PV+���/�͏N.�Ə�o4�OJ0Q{�W�	��/6��]�5�C�t����,V�2�x88�1B��0}��Y���z���P;������Kp�w�D�_v0g<���})��Gv`�YvXT�HL����u�#��$'"؊K���C������=� s��?�;U��Vّ�|���m�����{y�~<�k�S��b�*��f��-`
Y!\�gq!������F���BTID��Q\3j�;���Ⲫ>���߆0�7X풞[=�7ܴ��!�zRsF����_өw�V|��Y����Zʂ��D��Vg�N�yHM�g�ʡ�#޺czԪ���*tg��'�_)�pQ\C=��K� ;�zъB��j`D��R�^D:E7r�R-q��K�}a��ՋA��q��vV`�<3��ǩ ۷��I��G�����b�����q�17�]��a�p���qlVW��/ED�x�ڴC�p�sn���2���`85��g�p�6ᴏ4; ��[��C.�w�v�
��Y�QtQD�T6���@�2��Cy�@�e��$JGn���)~�ἕ�=���p㸭�Iq����M1��E��CGۄ����M�g���蝡\ ��5"�}i<�R�9��[�nHĂH}���1���{���FiYe��a�M�Nf�CꎓC#&b��z�&ܡ��šZ�'|I��6����L\�Yd>L@|v���x+��xN��Ɩ��}�kOW�h��d�> �׿�ϸ<�4��8�=�'�n�|���	$`/��z*v��m���#��O.��a�E$$R�v(X�#i~tz��Z_�8pF�I�e��D�N�#G��{9�Nת�\s�&߄S�<��r�R�����}�`Z<�nò�2]���#��|>԰;Z�哮�T�R!~ʭ�'��x�Yԧ?2Ɋ��8^o`(�,hz����ƾ��w�NsF���,�7q៖cS�Y{���� :qoٟ�4<���8�D>Б�U�Q�����H��:g^R������"����)�3�r�wԙ�k�/��0�����0̮���g#팱�-�I�#�A��E-�C��xp�F|z�r�IBv�t� n'-���pc��&knYӊ-���)�4)�
7KM ��,nE�]�|���@(2�&��hH��p��x�O,��;�v3�}���|�e�G����Yr��?��n�}�br���C&b����\�����\H�	Uz���ӿa{5X�T�1�玮<��N!��\�ђ���P�;d`��G�J�Kj{�c6N=��C��`�,g�����B����[�B�f]�ն1�̑�z���˶&2��Q��!K�������⛿$�\�0������8��Ń����P{���I<��|R�"��R�� �^�>��
��qgnT��a������[Q���l>�6�� }��u{�.Ζ��m76����kvJ�;(�QWzg8� �""�F=���云���^ZQ~"K�/��	���d@���
�QGX_^e�`#1�BL5��_�ho��M��d6k�z�J�	&��N�o��eƭ���$���i�'�t캊,�D[�� �V�:*�T)J��%�uR����sP��j��-d\���t涞 �2;ӏ�������9�����u�Vv�^� ��}��R��Ŷ�����"�|��g�;V�9�ȧ?�+�N�r(agL�ǘ�A�+cO�\�R�h�����6Em�������c�K ��Γ�7�LKY(E��z�9�%�]~��G��j�w۫X���k嵺xc\\U���ى�����z��P�c��)b2�N�Z�zN�-u2��A�m�|���Mn�݈[��1����r� ������$���MFOꒄI���U��+NS�,0��N�ER�s<��4�5���G�)__�E�	C�>4(��e�!(�_�O�7�DG��$��>���|$4.�q�=�^�w�Wl��j�$���	�9�?xUk)�8�t���0Z��BwN����'�P�GOuc#vvۅB�M2���I���D�1����%qv�-$�&��ӝ�9�?�I�N{n�U��3T���ǈ?�&>^�d�En&�Ϗ�c�Fd	#k���덴Y�w.��A_m5C?�%@8U(ϐ�c%%:���ٰr<���9{�ЪSF���)6���<C�PΫ59�3��w�b�f",8�	�k�ǉ_�
#k�CaӤ�c�&�GP�{C%����������ڔ���쉚�ĦgR
�̽���h����P�7��a�,X��/f��'w(,�Q�_�
B�	����v���MY�j䘙�_�``��N$�Ig�2m�ǖ�@�B�)��|z%K}��70�?���H����9P^��zI��І#����{�#v���vE+���R�8z��sxff,\�dco��z9򧐷k7�&������Z�N�JWK���?�y����4���8�HC琚FԫD|3el����d`Ѫ��1���tw������R�����l��*�s��]L��� �'c�� ��y|M�%��B�Zߢ,w��%'�à\��߶%}�O*7H�J^_~� �@�x�^eɗB�	j ���A������{�{yn��L,N�X����F�{M�%$�k%\��kx��9��<[�>��5�8OW�,��k�cyܥ�տ�*i�����w�۷Ǟ���pO��G��DR6ז�~�����Jl����5t�"h�����=g�1�Ỳ��$�.�����WYMm��]�n{��_�ǅR��?��,Q_GbL��JO����]�+n���V]�L��r_����b�ŕ<f� ,!�dǏ<t'uV���ڡo1�ߕ8��ё���L����Żk'^�*����m�߾*D�c�3�
x1y8L�M��MH �E�=�l)Q�ż�Q��R�b�vL��(Y�d����7�T#֒:�h����9�8�[.*98ir,am
��4U)r�)1`�"HL�u���[k�K���%���w����o������Ff���,���ʻ��{�Pu*�d/��g_�n��@ه[�;��,�gC��K��"��Y�U�vu9F�ʵ�~t�4/��K�B!z�_i5/T�(�������U�G���(<[hÙ|�fw����Fh<ϿGv�]u�����Q3F���cЊ�������P~j4w�:�;`k1� �	��'�WY������(��C��n��f��t+�3����J�0��(,��C�rSe���s��.NV�/�/tU�>�P����禱�~ݱ�"�� Z��s�;�۰�f�|s�]����"�i=�J��5��@+�h���%�Z���ۦ:��}hPА��w��K%rj��,��2�(vjLzό�޶Z�lv_1�}�g���Yf����yߔ�6�Wt���!y��0*p�DV��w<��-�;�C�y��!�=;��4�䭞���&j�g�smޗ�r�zA���ףծ�BV��y��}�+r�l�9�ס����&2	2��*�;J7|ОJ�^�题�)�Ņ�����f�75�D�S��J��#��i\��8<o��0vO�b��D��a95d*Mj���Q8���/	ur2pm���o���;����bZq�K�Oʕ2�v
�;�}z��;y��@D#����z('����s�|��`��IR��z�k�m*��lTb����c^�?���K5�G����Q#��M���k�,�Ctt�0����K_�vTX��y-~�n uT��(Oȓ%Cn���{`�w�|HU�O�>�>�������l�uޑ���R�!ڤ�
�p[�*̋a�y��0���I**q	����ݪ�B��>]��J�Y&�\?̯��8x��ޫ���jH�Jcǳ���S��w���\t�%��Xv���	ؤ�Zk���h�� ��n��B�y-�l��G�R��fUH.�+���J:,�=�2A3��Q�y�Dag��;�a#	f��B�kn9�[L�fܝHڮ��6�Rn\����=����^]N��ON�z�	(���R�֚�x��>���m�� j��р�_:�����|ܹw�zTw��`d��٥�[�[�}p��bo�r�Ţ
A�� �_����+�{%��K�%I�>��z�'��>��H��L��vİ��O܀Y�]�� �]���d�~���A��uEԹI5�8o
ư�d3���@���X7̡F��!�s��3��#��[�h��p@����O$�"�zK�Y$�N&�A�%�[@�Pl*����1j�*V��ݿ�ݘ�b;�����;O�[�]�h�J�k������7�AT�:4b�uX%���<�,:�r����_���u��Ц.���+�ѳ��lq�T/��=����ߌ�꬚y�rȲ^�+�@�kUm;1;�?��4�
�G=�/Ub���i�I\�7��� �mx�
�O>Li}�A7Y�֕���V�z��x��.��$1i@J��#�S#�!�Ϳ�J�=����̹iJ҉e$�SI��_Bޒ����Wc�M��-Y�������?� [N�.Eu��B���}����3�[vl�7�ߞ���q��/��foVJ��q�|Up/�'�& ��nO�����{���2RF������\g���C�uB�����M�3���>3�|/��O�A˃��������B�>!������l��YA/f6�{�3t�k}P�}��x�n�G�/Șo�~�%�@���叇#lw����]��|�'�]�ln����p6�����a�3���,���8-�t������!�"���@TQ����Ԩ���uL���9R\D
�(i�ǣ�ܟj���Co�5ҁ��!,��l��������:���m�$�����v�r�,��������V+�hu����5�a�WY��&=ۖ!\����3��`�f�jX�Ϳ��9��w��H�T0�'9��*u�JX�z�^�����<��eХ�٫�مg�A���&x�4K�A�Ӽ�I��N%ۿ/��ĆS� �i��l�9=��
��gT\$��,m�G>����Li�Ù���՜hL�O���V�E~l�1�}�� _�i�B!�/��M�Ԇ'
�4�3�x]��C�evڲgdY8/MኞNu���f;7��d�k,%Ql��	����ӐA��ܲ�ё��4
����p:jQ���\=߼�c�8�q�Z\��	�;v�f��؀=W*ms�"�Z~�s�Uםro��*���1aeC���X�� ��E���&��sl�o|.�D�ʌi�5���v0�7�ϻ,�����.^�XyG�i�g?Ix�]�5��R�\<�:��ԃ��Z!�
\"|a�6TB��>�u..����|�,bS��A%�Zc>~`�.�j!�p0En��_�j�����,�:�w�w}�M�S}�D"�8�g2�	f��0Mz�T�s����b ��䫅��'f�?��
ِ�O�S3�Gm7��W��ߩ�� �G�O���dn�2�́ATF�W��ZחwH6y@���L�FUp�$�?K�~W6p ����P\SM����v�՜x[:��L-��8�2PW[���D˼(3���S�:� �3�R�y�l�9����1�����l����Jw}�ne�mS��	b��0Ŝ��܀D�.��T��w��c�,R#ng�VI37=��Dzi�gtʦ�`��$(���D���Q����A��68��i��-���9*ĵ_�ݩ�	~.�D���<`��A<�Z�[ً����S�{g�&~�c�Me��w��Fv>� a��7�4@lIi\\ ���X�SV��Ͷ�zN٣���,�̄6@��=e<ZVW�YF:%�AT��9�i�(�g�z$Fa�*M�qP{�\�@�$�j#��ô�oN>��IO��sk~,T샴?P���Z��k`<S��Yo�G����b�S�Yئ6MZ+�0=7���J�GYĹ���]g�y�
X��Vվ�]�4��j����m�t3����01(��|�~��d> ş�0�dp�;�OU��17�ă_��`���(��~���kμ��Ac)E�y�x�.}G?s�:-SEQ�`�_������Vө��Z���te������̝=�͋���8�����]����W�u{�ƻV����G����%f����2l��}�#ΣVbv9�󵈋;.�l9���E������%9NگC,:T���7�d^�w���k�*ͺ�#�5�����>�oLd��c4�'�՟J��D��|�$��4����̌V���+�F�B�4��q{�o���g���5悃ˋǩA�	�Dq���aF����b-c�b��/ʿ�p��g<J�\őe�9�C,���Kf#�������׎��d�h���E���suIh�X��|�pUlqqr�@�Y�A5��ʡ���T��I��{b��lC�S��m���g���.�c
�J�\�85�f�����q�h�iz
����]���L�W��/ҽ�ĘUsjN3�	 �E�j��v��ǲ�ҩ�-z����|�11n1�g?22���T�?j0�&!���L�fF
��8:���F$Y��������t�����੠���C�ړ1J�?���7=���Ό�L���9�$�"J�}ת��QD���ʻ8X��+���n�TW�r���0����:Cݺ�������P6F�hr�DU}Ԏ��b��k�Y�Z�*۟�r/A����}�	��[���c-���
7p �%+�aE:Ψi�_�s�I�r-��
h|�=�B�r,WƏ]d:5�8�����w׾�y����7r�����:�\�-�0�)��$��K����j�����<�)�t��<����<��y�M��Z� ���$���?I:bĚ~����^����.[��'�sq��=#�o�r�V|UV�ڤl-k���G�V�_�f�D�q���j�+W�蠮z��l=!&��L��@�?Q?��C�9K�����s��L����Y����<�Ǩ�wF���\y�f�(M媂՚K�B��3@�(=K�Ҝ���S��w�R"���uY���Aa��8�8�����*�a�d@+q����%lR>�	��������� l@���3!�B.�]6�Ԯ��eI3R�p���ޒޭ���  �9�x\N�H��x=�)�Hn��o����lc��u45C,���&��~��cqXw�z�zQ7h%�
��w�@C�Xo����7�~�C)y���Zq�]0�k�	l���������zN���Z�''��4r�$�\V�C�6���'����t��N'?���Y�+���C�ٌy'@�(�`�]����n�����$+T�`/PG���c��u9ca�^[CCc�0^�σ��韽X#�>c$c�Ȑ.�r�{u��c���b���|�ujTqMmMnELe:�@��p����i(Ԑ�9-�t��>YG�IJ*y�� ����K��"�6�(���!�IJn$�o����|�e��o]��ܟU>Hh����#�o9����g����un�vs�	i���C�i]���d��]�r�,v��~`f������u����G��|���
?'��k�=��������)�bHTI�. _OC�6E����Z뫵���4���}�,P=b�e�=:b��y* ��8�n�Щ3���s����x����yl��4������7_I 	[�2�����:mv����o|rm�����w�
�������Lv�c����	J�o��w.�)�w�=�5���Kk� )B�}�g������3Dw����
_��D5�q�)X q��H�َ؎z�2a�Ҍ����?�'��Scm��
�i��`�V)���}�lfOc�&$�5��a?e�h��!L+��MĿ7J���׻��ݐ�G�L=��2b��_���8��(9e ��b���f��ׂC[��0�r������v�M�X?�t2$_�y�"� You����s�\4��\���榿��8�fe���"�(�W��<=������ml�io�zI�9E4�"�|�	{��M��Az��1}�1��5��mơl�jv>�}�K��#�q�N���])�6�����D�� ?�����������=���EG����]�VX�p���*#ti�C����ON�N�}�٪���t�؜�`m���:٤���1�N�LT��a݇�e��s�IO�>���aQ��pC�-�w݌��-VS[����~+x[R� P���lix�&ix֦ř�B%5�l������e��cG~����z	����w�+���R�?� &��@s;X�w�1���c�
:7k��t/Me��Y����{�t�RQ���4np#6��ȳj��QU��xޢʆ�[�oa�qE{���_�M�O�P.�u3i����'���}b{G����b��n���Q|91�^W���I�I�����ާ}Dë8�'Q�J���Rd%!!�$�t���+"�ݎ�&��f#c������LV�*C��9�X�O�9���3�!�w����l7�bGW��:�R���y`�)����Q�]��$?���5>
r�����M��TN/8��+�����N��-���l��a��X1p�e�^G2E�5���t��ިT翇�-dh�v�K]���A���{�iǚћ��ޜ�0��c���ۭ���^�~��9���W&sC�ӎ�X��j pl�k��� 4��AO/�i�&�y&@S���	��� �	8be-��w�'Lԃ���M�~���H߲W4r�l̍������:����{ai,݋-�m{#-D��V	=�2	�Bv���M�_����M[	sCA�T�D��a>��A��}}�yI>����γ�%���S҂�i��	�z	�X���ςM)N���G��>�g�=ۜ���^E�h�oj.8����>�2˒������E>.P�|Ssh']�}����1�u"8r�����ʬ4M�4痃lam�tV�;�[�9���6橡����<�9�0��{�lfe��;����<ԥ\�&a�/����8��Ⱦqg�'\1Ps��`��)Fl�0-��&��;�$АE;B��΅$B�TY���#L�hiM1v,w�v][�{ ���6�Ö�B6����BV�PʅK�ۼ��W�sBH�'|ָQ�u]?��e���P��o���MZM�c�Ӥ��W;��E�xg�WI����r������Ɋ��Q�Y���))N��M���	"YB4�hi=a���JJ����O*��~���t����z�)d;��X�s ap_�U�UwG9+8����2߰c4�opru��D5���E���"���	`��ky�"��<ݴ�&����+:����\��ؐ��g��)�X949�����ڼ�IF�mWw
����N?�4�M��v�b���t�N����_��֭��W(4�z-#@����}���Q�Pt[�%��zڃ�8%ϵ^f�h����&��|:	[v�G�F�}���XG&.lI�0�R\G�f�{�}2�_�߾}�Y�3b<$A�2�p��H8wXi�˄d�9���N�K�~,ϻ$�mw�Q���~h�ӣ���-���N
tƴ�_^��������?���^���U�y�r{2���=�a���r��qO8�|����� ���a����o�!����7�J���{ay�T���Š�||W����F����4r�2�)�{־����"姯��:+���!���~ E��-�-�7Yr�ʧ���F����%9�ϵ��Ɏl%�B�ٷVu�ƽ1]��T�$R�Ĉ��m;|�/o��>�4���T�	z�|��RXX(�#�i�ьF��t���B���"�k���`��۱��u!ҕƳ����FP,��?���ܫu���.���|��+eJӈ��&�A���v���,i>=�e������O���i�Em*�^�hMV!�%�4g>;�!�x�*s$�Fȓ��[ʁ�bq�K�������� �UQ~�a��\L�$����~лSM��)g�R�����y�H�BX
��3|%�!���x\P����(Y*Wr���#8�xУ�#GKvc,KvRH=�J����(���J7
/���v�'����M�p���Dyp�sI����V�gQT��H�¨���ԣ��y�[�/:�h����	o7ܾS
S׋��b-�t{fQJ�"��W]&%v=a�U�2�ý�e�,3)�C�i��A��]�0^6�M���*�]�E��������;ڽ6���]���r6v��{9���Xh@�>�5���Jb̕7 a���J?ͮ,�%ē{���Q%�x�!�x��?G��*����{�Y�^�ՖJ�XpBg��f���pa@�D��9��RB�KE�V/��D�!(tJ��nQ;��
s1 ����-�B��+��#�8�p��6�"F������aQ��7�#{i�R�G<�ixa��{T$Β��J��"��0쳔H���y�y-��E���!	f�?�9ԓ9�����3}���󯔍�G��P(����q,}�p�
I���9�n#�N�]TdO��_�z�v->z+�k̔�ofTl�da(�UƉ���Hwc6$T��g�R���t����T�����ow����ߦ�*,���\����{��!��r��p�^�,.
����R�bk��� @�WL���:��Ǹz�鐷�Q�:�����7&91~9l��v���Umm���M�~(�� I�V�-�#V��B��䥖<�'n� ����NA����m~�J�0B���p���`}zRUmq�M�s2~a��8rUT�r�/�c�T"���k�<�l�R�]���y=��23k�aYGo:ƾ�TT�s��Ė�Q�/H����iV3U�ᘘ�f���1nbbAo�A�� Gz������W[������#1�V�� �gٔu�e����I=����2fm��8
a5�4d�����6 mR)��_[�:4��<�qI:�o���Jlb��uk�k[��0�J��4%�����?@nM;u��x�%砩�M�p�.bu�q-GS�r��������D�g��i���f��^z5������3��O��\��yb���w_�;�Aٷ���ӓи��`T��A��}���G�$�&���u;ݿ:1Z��2�`�?$+��C�f�_�H��4�'�)��"2�b� 3��`:y��R���;p�Se��q~L��%qۆ���w�&L5�1'J��n�u?z��]RTV���7K��]z�Fg�IoyQM��'*���?����Rȏs��n��U:�>�x���*Y��ъr.��2��g/�Ύ"�Hl��e�Zp{��@!_��sP['kI���q"~�c�꽥;fLV���4Q	�S�.E�wq_՗��߀�R��qY���8z{p����kc�#��ԋ8�lF�d��Ǫ}�FW7�O��m����-$����7��U���I9(@=K�����܀�&�0n�����s��t޹'J�A`U���l$[��<^:��)2Ǐ���~�A,A遁��I��p⩈"��4[��F���g3M]>���H����sf��6.�%z0�`���y�'��"E�B|��� �����@���{�/�@59!u��_��)�C�y.y���zY�xO|e�����P��+��	E������Q��C���%ũGtU, 0w[^^^dd�?��Ӷ/�)�l/#L�".)iF��@�vۗ}Ƈ-M"U��p6��x�g�;���̻ھW���o�^�� ���e�T�8V���I<����vjy��,��~�e��ߤ�	��a	��6c�u~r�v��>��j���$Sm[��D�<�h:�hnwf�l����+u���k3q����a۝�r�E�8�� " ���+z#��y��}t��drP`���^ ��|���p�ij���a(����~
�s�f]$Zf»��R�a?Gbe�m������d9�mb�7:�`	1{�
���ge?�q��T�en�;6"����H��A�ڹ�E�a��O��6�6%-�Z�q���m�ʼ�����5h�8
�C!���6}�~~/�_�=^	�πږGo���cWBs��g�}x㚥bGw�p�{�kG�ϰ{����#%��&xiCG�QZR�o<�4p�z�߷�fPDs4}����\��p�}V���!�2��q&!������c�51a�{�^<��\P~)�;Z�\��T�;�7"��J$�����A'�uԚ���w��+������ ��T���Z�o��6k���V�m��a�.���Oe��*Gv(��m�;�NZ B{f�IL�M5
�K+���_CP��GYM/���Y���5�A�p��9�2���,C˕];H����sa��V;+��č5y�T�R2D<��9����Rֈ۳G{l�in�?��YYY`�J�(P�S<¾��������PFgE������p紉3���;gu%o�F��B� ѡ3�<�ٴ�f��iPم��]�#]���뱈.N��7L��uR�����?QH�͑g��faW0>��$M5N�����P��AQ�`��+��ΰ���s� ��]�}
������>�fFs+̮3��]�p&navz����|r��h��.��\����

�i��BLNګ�z�Zgf	ܰ��è�mѬ��6��&���rs{J�h�kT�9`��<3F��Y3��2����!��V`�;�T����2x��L��Q���f���ڴ�чn�!RN��w(K���`ܞ�%.�,�e���]�Ȥ֟i關q�_6��@��_���X�2���N��;�+f�S~Ȳ�E����g��؜<��sǐ�8�� �Q���i�Ii��	���)�U�4��(����-Va�7�yG���W����ĎS���<��Z�����j.��m<ߥX��O���d���.z0���չ��[���^~6��z	���Gm�s���V����6
.���Vd�@y�,\���g� 2�t�$�12��J��o�O_�7�4��\η�f!�6!�����c�6�u��^�Lgy�I3+(�	��P����-�Q��L
>�96�1K뼱AöEw2��L�\���t��A`��8�T0��PK�I������:�_bđ>�`�O�Wq�=Bhi�C����;i֨�"Lp�@Fn�q�P:��Z�����Uܬv���bw1�<��[�4��pFRLp�qd�G�y��ж�*��zH�ٺIn̚y3Q���i�֛�<ՏZ����p瀕�|j�B���1�z���8.��:n�Ȣ]߂yUX��ñ������l�u�[��61�j)����;�ST=����	;���w##sϬ,n.�/!���D3S�Ӎ�v��������$�4	�
��+bNG��D����+Z��a&�#�?2�.j�9��
5K���fA)�m��մ��b����O^�a�̈Ƨ�)����Ւ���أ\�͊�ݠ���L�}V/����R�����46�]i����%�;z ��(o��a�&\�И���hљPJ&�w^*<ĸ}�BRKKK!�����$���֗^7XY�rN���wY����Bحu�7 �!�w٠�t�K��.-Q���H3B�N�Qc�[��AD�0|�� ��F"�z-��£YL�5eE�É:�y8!|}iڻ����L�s�z�c�:Z���eAg擟v�޷u�����O_�v�}M)������w(P�X� ����
�X!�J��Z,�]��~���f��2�d��=��wם���`snڹ	�;�t�M���|G�pN�T<��U&QLY�Qn�2�9[�_v ���upበtC.���*��u����Ȗ̯X�B6��������V��\<v(�?|0�ܖ�r?emr�:����1��AR��8��ܩ���OVPo�Qg��~29��2�\!�l��	Pe�"�hn��у�ќ{q��稡;i�,�[�Y������+�� ���O����6z����Ӷ6�{�nٿ��K�gu�ӂ�?Q'~�N��3�"3�m'���o�t��(�b�!������ܑh�����^��5�6"���E-u�E�,c����+���P��3�f�����m��W+�$���M9�ݭ2.��T 5��>-V���|;=P/�l���(TG�Q3
�nl���E�6�Im�&H�!~��{�Dl���&~����(Gh�5���i�i��Lz�����%)W��q�k�C{��1mITkwjz���Ժ���̧�D�m�FmT���!g�6sMC!�DD��>�-��Ww8!�leVG�fLX�o��D%���+�C�o��p�LBJj|�ZX�AY����us���o�����צ�Ǯ`����_}E�����CGr촹.ς	���<��i
�kU1���x���1�����95y��@��7UF���N7g3 *w���C-crlX�گ�2��n������j�+Wz������qf����8����a���$$s�I;0��;ȶ�Cm	�+>��[�{���`o`�C�J��G�=?�+fd�[�T/Х��sݘ��ZʣV�f�5�*`&������ԴC6���p�A��2�hE�)l��@���3ؘ�ׄ�Y�~�_�_����U����M�Zsek���&w���:�/��N���x�bf>�Oʹ��^�+���?d�]p��=γ���)��-�ǫY��=�5��gf�Xҗ��Jzo���b�t�~=����I��]_%��!d�� �{�i.dF�%��E:w��;=I	�8�ngh���_��D��:#�k���@n�ū��;W�Z��΋)��3�Zm��[.�3^p��۾י|��~�ɣ�hQ��u��8�h��><��&�r:��{ؘ����JL��_�R�9�蟇��Os�"ȈOk#"Z�"�����	Z�H��]�N��#ve�Է���j1�-�.��6V����>(g�.��#�׀�$�Yi\j.��:	��Ϲ�[y�Q4�[���*9�{�(�Z�B3S&���H��b`B]U H��t�mL���B��Xt�T��'��UҒ7\0�5Gzb_	�dud���ך#��6i��	jQ��=�?��������R זOOG�������������l�����c�@���v�+��U���,�m:i�y���q)�#A���1��hɞ�w�Z�z���f��~u	D�m=���N'h��-ى��a����h�����=�P/Y�z�-+�T;Wv��)�g��,��]��
�#S���6h:B��zKwK�9��YGc��|�;��:&���9������!M��{́޽ő��c{${r�3ߧY$ۓ��sV[P�K��Sݖf�W=��Ô���6{V���m���O�*U��Z[r���e��%�Lzyd���r"W���.$8F��q�ٟ����K�wY�ҙ.O���x ��)��V[�/�>��wF�S�?ASV�*<�,�6���ӝ�^�9�;M�Kľvf����H������Iݹj�o��[�~�5l���u������u��mݛb���_���kFIU<�r1b�a�<`��4�����|��j�<U�VB�J8Ҽ�3�dH�U��h1�4F�zӥ���0��B I��!�h��@��6�H5Ԙ����->�*���,]����h_�u:�bu��f��}Tx�oJZ�&J'�{���ӱ��������2y���?�N���ԋV׭���#�Fj�@U���]�+a��\V���0��IɌ��$�ѳ>��@��
Nz�Nׄ��MY]�3%�ߴ�i·hA�fFFK�,�Dd���K7do1��?B�@�Ԏ��}Tx�<����`����f˟�dq!!���!7���\�X��q����3-��m��hA�Z~B�IaR�fR"ҋ2/��T?��)+�b�|����k�>��T;r���lv�B��/���`�����gk��
>��lg<e�Cr��D�V��5��E=��H;��Æ�ME,�%Ӯ�K�@�rmC,S��M��T��U���L���S�N'��㭗��&H?ܸbF�.עqz����nd�t����X�]˭.v���H ��
`1[��t-X��,p�R����K��mc�����h�(�����qZ�������_�0�@����t���rt>�LNL�f���Y����"�i�=��8怴��
�������A�Ԏ|�m�˦}���_� �X�Z���Pf����֦zi�qL=��6�<Bf�	#H��߸?(�����3VC#��~����W�S�4c�_���r��"l7c� w� �)���B��6]��B�O4bzi �4�^V��;90�~^nkb���2R�~%��b��r)��I	ڌ�os�J���M���G��d�/�T��RR�b$���
���e'�爼~��(��)&@��H��"�R�t3E.(��$�-^�&�f�����b׸��9��S�����OE�;�7��������dP��G^Wb��;>>lP]�U'	A�q����߰*�3,o7�C�ۗ��26�$�%��k�9I���?�a�2v�)}������}�������땀N���bG�}�
���`�A9���.D0)[� ���~)�X�/�&Y�s ?�~��+�X����$�)";*�#���lW��7�`�y�:i��U^I9,�S��<�ɒ�p�/^�Xb��'��ns|]jO�0&�$ ��eۖݻ��4���D:��� ����u�u���B�؏����\��^��%#Sdb��Zo#0�G"��k0>�Ƿ�,w��0���s��c����fסdpc�/"����\9�6_T	E���q��3�gU(k����"ϮV���YJZ���2sT�C�|��[�����x���xց�� A�!�y�����9��LFԚ$Kp6.�ޡ$����*y�)R�znIێ��;��ib��v�~�9^t���{�Os3��D�*�$��)#�T`���sF$.�#Z�zW�H����8	=ذ�)�_ �K�?�n���l���\s��r�.c)H��Rﲧa���^��2ig���'��f�ң����e'�;P�їd����v�_���Wv��+���6
�S��&�Q������?�4:P�ΑIEl�	����>X��վ������=��Y�4A/��63����3�*9��C���\�� D �#8f$����
��޵w��\�ztG�)�e ���f�M�P<]*���:���8���m��̊�o��O����1�K��O�q-��i��#U��S����p!���_�Ut�/����̍�"h��!������}p��}�b�Z��'���d)��@��n<3
�~̟�3�ʲ�j}��Uo:�[6�����l��6�O����vB���H!�w�5��s�΃@���.��!t��ￃ<;0��l՝*Wt�S7u|�1�:l.�́axd#�ɢ�&�c�{��?����7�6`V��㚑�����o��8V��q6�W?`��eWd���P���꛺Q�Oħ�����q�0�� T�k�8��{xMk`�@3H������C��ͷ�}���
��-"����CJX����R��X��n����?��mo�b��8��#k+ip~~����}��K�a�QE�s>!�<A��*�_�F�{S��N�9�x��ÿ��s�4��rp/ԙ	ˎ����Zj+�i�Z�����ڒbJb��\&ݜ���X:��agG�E=ݗ���z��f<��~�I���mc~�"��������ZIh��%�w�zp�_�>t��K�����A��۪��T7���ʹ@�������cF�nݥ��d�^%�I�K�l^�|��D��d�U�BZ��:�|�[w�A���Y"�q�H�5Kr�����t2���c���pQ�2_��n�턘7#ݶruu(��v�ǉ����o_P����%��D���:n�8�p_2(k*��w\�I��_E��A' �矛D�:y����+b9��[�gLFG�U�4S���!�n��M���A�SY�����KǚO?���ki`���s���Xg�@C�������8��Up)E�ӵrhp�J9A�4�����_t��6�M+{'{����o���&Ã����6;�X���5��I
�c����ik/�ȓXdY��I����8���Cz����� ~�Ҽ�Q�N6��j(�D�~ن�4��Ґ7_O�/��{��ap��\-v�=4ۚ4��Z%�}�`Jw�����\�W�s~��S�frٌ=��Zn��q��.���6���b���QRn�?�p��>�0n�����bj�q~�
S��^1���l=��D`s�����&x7�%ν.�
���4y|N~!��4�� ��M��QeoQ�p~�{Alk���	�MX 1��v��`���H>�G������yԅA��zgpu�b!��b��22Ys�.q,LH	��@��QG�0E�Pt^�ӵ�k�=DN�,��T���恑���T�z7�~�}F"EP!.�O2��TƕHW7k����1-�c���~W�A��N]�;w<A3�	$�)�
 H����#�1��������bR���~33�4C7)��}[��_.. ,�D�^@� n������'�<�u�������߮^�$7U�Ys���ϐ��3�[���=�i6=������l�F��)BPWZ���~)�����?l��%�4�|�V�I o�9ߢV���b�
��i��3J5�^���KZy����HV@����-n��3��q�p�±����7g�CW�ޔ5J�Dg?�o�7ۤ�_����.(�����Oګ��K�a@F�+b�tI��L�z�G'��i#4�xkύ�E�R�ã�N5y]VG��J�N��S�_ ���a���7a�*΋3C��,J�ښR,�s�y�]@0��o��_�G��Tp�:���3����׾�&���[�wr�T�: ���-��S��_c�1�ҷ�o�<h����+�9�Q�r�PP�B�9���S&�ﻚ�&cr�-��O@K遬��j9O�=[?�j��	���q���3�eTgk�Ii�kl7��hg�q)~�y4�����i7�HS$4&_�C}�����F�w�*Vș9�e��{Z��V�������^g�%��i�&�Ǣ\��s�E����������%'�gsJ�5�/��z������5&aIQ1���>�5UP_݈Wj���o������r�	��t~������Ҽ���c^��b.�GU)�$�͛Sa�r7(�K�n[���'s�o�_�w�F�L�`������h���V%�!���y��?�I"�\,���{T��Rz9�V��o�-��q��t=��&��jm��k���&�H�<۷Mt�lA�q`����y���p����\�z���3����\������l���w�Ŕ{�RtmBV�ƾ���k�ə���:P�2�A�~J:j}_��d�;��������>�'�A �h�bss�q	�~�2k���2���]��3W[�n��<��z/���0�d1a���|h�]ck�o���y��-�K��`������&�J0�
�5!T#�)��9y��N��ɭC�dHs𻥩'�GL�Jc�����ip��cB�\(��#q#�mi��J!�qԻ�hW������U�0C��o�N�����y�o��O4�},ú>�d�Ȃ���z�yQ��L�<9��oK]>j9o"�rm����EJ�O�ޝ11����oe�����`u�OaBY��us���văl^�1a,
�<h��k���y|yDA~���%�ON��n:�ݵ+��mܨ��|fȃ�K�s���f�֘N�MY��%]$!W�?,BÜ���z+�feMm=��)z���?W�%<X߭�����%���gCC��;�wT�ؾl.0��P��k+<�l�PY����P� ��Z�G�7I�<�[�:�`�t���5c�}�4c?U������2���sD���㕪�[�QC}ݨ�3�G^R{��ͫ���r�֗�X?2���[�#8��M�뉞ku�k�wܑT�Ft�]��vmJ>~�J
v��^�<Y�IԄև�̪�H���ɟ��ƫt<6�����5ײe����3A0PW�F�Ҝ��2�^Dq)Tt����eI�X�(#g@<�m���QR11m[�N>�7�BJ��n�"E��T<m��c���S�Qb9`����O��LM�I��I�A���0�Q�����i�/��k{��2j������6X�Et)�kW|a�Ý�������{�ڔ2B����#���N�8Bv�n (�i�_�����Q2ޟgq��HB����պ��'dD��U���'c䃙�a�=��򺅘sª�2ƌ�M��h��Q�s�Q���-��:#���sE�����q��O%.�Y֧~l��1�0�#=���WD�{�v�::�m�>:*�sIm�&%�!��-�%��YN�!�t�����H�mWTeqr4[�K�Rq���WL�=x�VV�6	t4����n
��[l��Fv8z�Q�?���5�M_�=���%�Wr��҆k����#�l�(�Y	.�ӷ��1`!���b�H/��e�m��/%��֧>���L��E?�W�,ζ��7�BS]�4L8�Xtٚ�,,�T6�q>`�w�n�HB�����ș�/]��[��w=�-�~N��ri�#o��q�]�e���E>��(�<���^��c|��k��w!ۿ��;T��s:i���5i�l�/���ɺ��u,�xu-����<M�2�z�ɏ�%��Y��7�P%�>�ӑ��B[U��9�����`V�3s�$s�o���w#�$䣐�,�׻6��Y'\!� ϊO�-���y>��w�U���G�D��[]�_RK
�)�ӥf�f�FP�,�?���6��x,�܈ <��&4�E�k7��jx�.k�@�&��#����ՙ<&M-��w�cK�>�3Y����`w�6C>}�a����ugv�.`����P��w}�)�˃O�Bv�tͬ��������_�ɺ'����A�:��o�y��NeE���T݀�S5X��ƻ����iƾfu~�@�����<u������2IKK��_���{mB{�6��x���~��k�
�� ��5�.<r;=��&��:Y��9��I�x����CnR+E�m�61���������%��\�v�������U1s� P���8U�[��q������~/�������Njdo�g��8<��SB�r���{��@[���� ����?���j�X�i��z�kt�_������
���teC�#[�7S���1��O�|�S&x1jm�c�yZ������Q��B�3 G�OA;�����X�$�hJ����T� �z�V&��9���Q8&��1�:P�p���Z�<v��t>�7��]ko�'�RjBi�u<�E����l���
٦B�Ts
���^=�=jM��v�����;zbd+�lJ]����s~�I��~.V�k��+�Ԛ�l7�\3����.c�<�9���0x���qŜ�����x:/�r+���%y�.���ￕ&�R�ؒrr��,,�QѨںڒZ|���U���c<�ؚ���З8�^�e�[��p�Ѷ���5fE�e�����卜N!3�t!vQ�`pW �֏����S�,��Ʌ%������h�KK�_h�R1�ejVo�<O���t߹\/yX�M���loE[�s����R:�n2�5����
�Ey*�.3=��y��Yjj��diT�[��"pQ��3���6�z��T^�RG�E&��d��N�V���j�è�Jo���bs� 1�7~��7�ـ�69N2��n}�ʠP�H$/�ī���ɽ�h9<P��n|���ooK�V���	Yuݹ�V�o��LE� e0n�7�18�k�*Gp�t��PA>?\y���m�9�Fl㑗�C)���q��"2t��Xb���i�=|ﶶə�P��#I�I*81������N�����}��F29�t�W �bb6�vr�>o��> /�j����!݇���]�].�HBw?{�.�^����0�?�9������Zym\�ڳ�0A��+�hȠk�����j���M<�[l�i� �G�<ې� ��_	���xT5��H�X������0؅)��}I%�yGKK��T���/�R��,)f��1�e�r|f���L�IC.~I�$k��O�����rG�����$D-���B�h(�Dml������R�=X�eqab=���[z���n���}��pX�+~��x��������j'/D�q��R��7f��M��)���G��f�g�s�ޅ���=۷}��G�	}_~��`��BZ����t��,?v�ɷ1`BR�.Nsg�˘r� )����~����3}��_տ�vj�E��Vw�и�^�z��FI��:�0zO�,�z"u���hn$�ĿQ ��cQ�+a[[������}�[J����H������р�c���{�ِy�3�����L����`٢���I��)�ZѶ-z��o����^����ң��·
��Dc�e�TD��j�Q-��H-�؏��j����Qo@u���'W��D�k��Pj�R԰�������a����(�C��Ad��w���j��xQH�U��RDj��*@�\J�tn�}2fD���WXI���+�>^K8��9Ҙ�5̫bb�@dK�%���A��I{��!�h��8��ډd|�dۉ�%����$H�nԵ6Y���m:k�:r������ى`��s~�Dy�W*2�Y��U?"C�B����+m!Q��nnn���b�w�e��Eߛ��[���ܽ���	D|9=$6���~�������+OG{3a6�9 �ؿ�s���<�:���1yvs۠�䁈a1�4�����a0Tb+�D��	·� ģ���}U�#����éA���r؄�O´Ԥ\]y^:�v��r�py_k3IK&��E���:V"߁f:�%���z�LD�Uj&M���6�>���f�k��nsU�Ƭ��Y�� y�@�#������%֣*��6�vB�����N�֚�+��������9��� �F�-P�� �@O�0��ӓ��Cqa��H�A�ȄM�]�E�RO��[>��k�R���f�Z5<��p��B4T��IH<`Pe��{G �vDX�jwEA~��{�ܑ�J_u�;���0X2�>��X��D(^A^(�ݩ��闫FF���Y�M��x��?�~��	łY�kD"���y钥Jl��\���)B
LG2��)��'0^��j�x�G8P��Ҧ}28v����1�{A����IFJ�T���@BBZ۹�^���4���� ���p"ŵ� -��T����!����~�>|47UI,�m	�C����|���$� G�m���>��;��XF��S*�������&�У��� ������]���!�?����EoVC<w�<Z��5���ns/��г�����*+��{TM���K�+�z&�����'h�l���:����&���_u�1;���2����Q�}2�@C5@瞴���k쨨���),�C��:�~qqaz2��;��� ԙ546Z�}%��m����mhj2�.Q�m��5���@��c�0R�+$�W�� 2ۏ��oн ���`�\��|9�BOW�t�m�ԭ�EG|�jʔ
�X�M+�� ����f���^�ڬ�e��W���L�+��XR��zH�h�=�'5c�{9�����A��[���E{
9�"8�a�/���.�̨�*�؏f���H��,,���=:)�:��KR�̩+��]7�SVs�5ɬ�����W���;�Oe�#M���W�-��k���BLPo9��{Y'Xq��8K�;�-��pZ[O��8�^�����-�|����	ψ���H�~�ֿ�ϙ_���!�r�{�6 eˁ�0`�I�к!������թl�h��������3�5���+�����s�������Q7Sm/U}y��t�Q��UPh��[b}�u�����w[e✝wTj�"��Gߢ--K�9^K�V{O{�C�>/C%���v&A��.�R�$ta�a.��Xr���
j�Z"����(�j�������k���i��֥*Z[[[/G��X��CD	�~u(��s},��*a͚��G$L�7��Ԃ[�l>;g(`��bw����֔����y,r`����1���\����y���<�ix��M����+��nŮ��d����Y��+����ى!�h>�Ǽ.���@�]��g|NN�K��"�UTa�6�AhE��
#�hDe #K��}G�t5d�}���R��[�Q݁����G�1c(a$l�9�ts1/�����l�[��||w^�'����p���p((�]��,x, �99�hk"}�U'@����t��&(�E���ϖ��88��uk2.Կ��:,baa��:���� R]����"�����Q���n:� �t"ZՉt�'C2ЇP��ֶ�8�G!��R��lmp[O��� ������o݃i�A��:{�6��cҤ������P���nӐ|۽��Rot; �*�@I��Ҥ��!ߓ�j4�o5vKQYd�M��,W��ӓD]E�7���}�-�����#b.��g�4�).�M��:�FB�D���±�Q������6��ѳ`q�QPJ'�~~J�{�=��3�b"�=nLs���<8.i)�DO�9� ݎ
er�]>��[�,�B��#��o�[.w��;�����$�ߟ�f��E5�a�G�-�m���)��~����}?�|IWz$j={�_VZ��Z9����N��5o>���@��]&��6q�%$�;��vt�uIc���d��0��cg�x�#�|����mh���z�bd�Uo�F&����,�LČ�P�`k5���SmG���ҟ՝Phjz:��d�/���0����t$�����KY{049��_aޒ�'�'�xOw4��Ki������`����r iU�&�+G1W����U����� �+�e�܋���cQ	��Hb���.wG8�?�­5D.[�b�B���s��Ė�Ի����W�W��@퀖zk��N٠�o_(��g�(��g�{�3��A�6,��8V�8DA�\
��G���]<�]����	�p�\A�f��~������^����;��@��Zw@,Byhd����nt]	�IrugN��tS`C�x��gY��2,cbz�u�����ܳ�yKI�:x8�vg��V���'79�B(6�XI^upu�Ĩ Гk���>X`Bp��C�2�Á���K��5�����D]2�RM��u�J��<�1�f�aw�� �S���kg�'`_�nu&��e)�/�U���GH�iao�!-�&��_��)���h�q#��BgCl�	��
��@r<zy���Ef{L����ME�Ҹq�K�,�䞣w��]F^E�(�U�b�𤋮���Í`��`�����|��������&Я��0c��2��3����}*n���K���[��x��WРұ_4O@#��ӊz��S^�5 P�j��CD3=�;Cz���*�xߪVM4P���np�Bq��O�u��)/�)OT�f|�@�R���-Jv=�v#d�pW�� � %?/�VA�u�.����&�$�`��#D3�P��t��㊄��B�1�����́�K����y����/AaYș8;�<��[C���{|�uύ���x����l��r./��H.2�$M^���}�Ŝj��ٶ}�IYv�E:k7ϳ?⒱�)�id�~�������/���lm��`
z������q�} ��8���u�Y�o,}"4AU��*��Yn��,6��^ɩY"�^D�3�Q7W߄.���9.J��Fs6~��:j����UV���V���[+��ot��m:�W��M��<�E띉�b/�I�S;#�J�� ��\�B�<'�A�ir��Na�����煉l�K���ިפ`Ѓ�U%BvE���`,�8n�W��#
߻�RO��)��H���y���ђ]Z�t����n-��w��)2��W?��A��'����^�Df�����vh���P��K��λf`wЉ0ܵ�
�=Rts��2a�r�g6�ϓ5AB���6��N�	b��B����r�n����/7NMvH�@&}�lL_���(�
�v�-��2���L���]5̿bDV�]�_Q��с^Ŗ%X�	91J,I����Ә��_Ϳ,�X��*�![P鉒�t<���gy���|��Y�s���(a2jh���9( ������M]4A��B��s GuǗe$�~��ٟ����#�.��c�$Q�O��"��:e��ۍ��;�M'���+�+�wگ�yZ���&�|��X8�_䉼~��ް�v��xTn�3�[9hq6�̇��r���� '��X��I�L���W�!�SDJ?ck�	mS��\�r�[�z���(���eu����AFLr���k���[X=�q�0ø�c��H^�v3=^��<hĘ"*A����Y��_4��%y�)���L�*�q�m��}�n�+\�F�����Յ�|Y�k�(��n"�Q�Au'E�)�$ "w[W%�8u�����Xf������LIG�WM�/�#'Q�ۊ��)D�� ��\|�7�T�߬����r���L��>�,y�m�Bs���Z�L>k~l���oL݆�6�@�9�~���Bd�gu�q�l�c:���3�j�m�c�ms�QLKo�����'��&鹫��O��"�u��W7�ޒ
�3!��U����`P����$(�ԉx�򡨵
�mvN��:��͸;��~�~��@��W`���t��W
��.���E� �
&��G�������:���vG��u�U��P!Q�ޤ1M)!(��@���Ӱi�>Z����D|�_�Uݵ1�2���і5�&����]�}�+>�.ح9���:��N+�Ԍ����x����p���ʐE�7������P|�8;�\�=���0����	���Y�������3P��VÞN�k�N��K���F�W!zЈ��:8`U>^����|��9913�e���~t��%���R��J�|�] �u�P��ر{�������� �����C�in}mG��������y���/R�2�_��>},+���Q_�#������N���j���h�[LbI;����݃2�u�4Jo�nsʜϭ���ytk��q��g����7p�xU�,k�%'����R�%(^nJKy�	4�1}Y|HZ)WM����n����@.]Q�"2��Դ����=:�LI
�����^!z�~R�̟"V|���U�.grwv��8,X����?����ִN���[���$ʒ�H�yR׽�`53�����5�p�ӓ|7�s��z�m�����i��p�`�g�U�|Q��0�8�@�c'�F�o5����pWӑ?'��]hO�Tg�����1Ϯ?���0��޴~7�h|q[s����m'�p9�l|������k6fV�3����h�A�T�&)���`�	��f�ۣ��$�IcL����:0ȷ[e�Ź����0A� l٘;W���n� F���]Ȋ+�����<��v��Xw�R�J��SB��	R�s@K�]��'�~�T�H���]�Ϣv�d-C�.��j����j��k���}�_��Ү`G� dac!:��XTB�?�ţ�Uh3��9N�5D��=&��/������-}<�5�Zc<��9�*)a�v�_gQ�쁩�ǁ�#���icJ����$�"o~�����~=��̡����!<`cv`�z��?��"�X_U61^:��w/5�:��y��֊���tл�z��朊#oo�ɖ��86�\��0���V��C�wF޵С�D������yk52���:�����*��1	bB�S"h����zI�P[iO�����E�D���/(a���w��Ƭ�g��tl�Ӎ����Y���ϑzH:W��6T\}	"�Y_PR�����)�g{����AtA���U[W׼?ՖHScW������xU�.�	�<o���
I�ֈ��**��t�~-��8ώ�
���� ��Wf�c��n�4=��"���*XF�u����[�$����~��\j��!j���TLd���(��R2���΂�~��ɉX	�t1[_'�^(�P�M�Dރn�)܁�{�Cz���`�$Cm-��TW\�8�z�16��!�Ђ��Qv앸��"�W��,nn˝�A	��OClՌ6���XȺ�=4�q��x�i��ZΈ���:-���(H|}�*K��l�a؄��1�((�-e�~�7���%�	�:����@�Tc���8h�7���E�lXz�
���r�Y�8f��+1��n�O�$2D��~� �|�/��p��K�CJ21_�1����rs��^q
��Pj;����j`�_��닉�E�G�i%
hd�uƐ�	��H��蹜����-���Ⱦ���Ͻ�jW/�}��oNܙ3�N�7�ĥ�$o�,o>\>E2���[�Aq�0$3��Ǒ��1WZt�I̋�3K��|�>6]>��=���Cw��&^���ZT��?�H��Y"����S����]�7Jns�+��C�-�6A�'��FF��%�f�ݏÐ��P����W;T%���B4�:���Eo�'�_�?�.还��~����r�1(���ɻ?='�����dm�;���U�lY[�����m�?	1��G6~��*z��o�[�}���pq376��1Ŗ�ª����"��!M
X�E~D���Z�e)�y//j��/ו�i�U��ݲ�jH�Ռn����P8��M��ʪ����'�כ1��*1���A��=�4ڦ2���j�F�}02�7_g���u�����ii>(�rO���0�)ҽ����9�&k�fub�ڠ�8H���ᜅ�,���Аt���5����A�JNx4�J����)��r���Y1]���va���Fp��A�<	))ࠪy�A�6JG����w� ����rl�MlUVxx|�)]_p�?�U���!}���W�]~R���@�7a>�T;_zQ�Y�2��.�?�_��������Ø��z�&q/p��M�Z�h���tTP&0`�q�n�9�.|���� �:P�$�N9n:>���`v��0�W��B��Q�[Z�y�
k��y!Wf}u���8�馉s�
� } 1��ݽ=)y�c���"����EL�Z|�,XP.7~�Gy�q�gu9s���u���7#����H�-^�O�������s8�o��$��!f5��qyh,��a���W0�+��M��R���I���K���T��ddrKKb6���CE"i-�]B�0�4�B�/4�{,�E�P(��O�X�Y���Gya�	�U�nK�c��ۇ���,���I��ek��Զ���+�E�'�$$�G�����|��8���7�W���9�,�hi�䷥qh�HnӪWgs�>6,�ik��[d�,�cHNC�rG��z4�DTa���OX�S_(
j+��"=<]UD3K6��{�ַ�?ؘ���Uڃ<$b�2|�-"�6;��,�KW}#��C$�Ϋ[�0F���q��P���-'�{�)�NA�yE&ވ�V�b
��)���6��R�6t�<Utii�����Z�t�!�O��{��ق�����&c"����Z.t_8������aV7�GS�(��,fTo@<�l�Qz���K�����:�f�S�ӛ��jE����հ��1�㎈
�|� {�m2��,Q��4�H�0���xi��+�f��1cϣ,�GU�uڼ��� -�F�;<�I���7���v��Q�/�Tک堫٦î��#�q� CA,1�~�B����%�a�>����؍ ����'yT�[A��"p=���ewW�r+�I�6TR�
)Z'+���b�����K��q�8�
K,8�t�V�A>�wz:J��	�82�r��q��m_#hҙOA�����;��k�d��F�[8���
��޶����>)x� 3�]��ǿ���>�>�S	v������LN�П9�aV�	����:�̃`�%FW����4AGG����aO6��r�	$aџ��}۷h��NR:˵Qk+T������ފ�u����c�T�Z��Qt�0ij�l�w2vv�e�WėY¹�)��H������i� �3s����Hc��f9>�#
���A��/�L2�C���q,L�);�c̉����@GC;�E�����j,�����M7eU������6��}�m>�z�r ٛ��[�E1�a&<�?��:*�����S:��S�.I��隡�SD�AA��ia�!��!���{���5���ଳ�����s,���·�ArA�7A�?ҏ��k��F�X��T����'d�Þ��n����]]</SLL��Ŭ�$��o�&����i���[Wv�"�Q�d=K�
 ���/݂�1�ۼ:|[ǥ��W�v2u����u9Y��u���w=�vࡪ�W?^EU���'Yk-��\]��sw�Z�x�|�@�����;{Z':R��~?$?�JKKN����P�@u�޼+���k7b���#�h���OMV��g���}�viݧQ���@1Gl�0���-��ڮ���L�&;	_��p�nl?Y��-�]��/Fŗ�������s��OKio�U�;��Z}8�k�gn�ך~���DZ�h���j��*EHb

�u4I�c�&��׳�lmK]��gA|�+��BGG�ւ=r�9�GE������3;4E�f�ŕ��ۿ����1�ϑ��$����������_
!��&���Fh�Pq�R)�l0���Z�u�⽞pu��x 	UaN�ñ�WN�$rZN�:V��y �p�!�ig!�0���G��*���Δ�јe�ϞKp�͇/I�d�c;��	bEU��R{�C�kB5�Zx�Z:��ӌ��v�������-��.�V�B����"�u��9>a�zZl��{:�-��F��Ġ==���.������]�YI�?�����Djk�>'�@/��ʂ	v��/�����X��U
���;��I�0Zt6�}��w-�dq0���m���/�ϛ}ha�4sE�Eg���V_.$�4٦��_��*1[�=�o�Q��>���c��P.W����yj�2�NVv���b���Y�W�/"E<���L��&4p�w���|�L�Th=��!��C<�@ ?��4I)�i�r@�Ԋm�}��{��� ��f1 �d�$D�~����H�?&���,�$����Í�d4ùJ� #��-��E�?JNK�Wd�s�G!��ݫY�[ſ�Ԛ�����fP�LS�D|�}M/r*�Z�uw���v��X�ť�njW�Ly�Z̨����¸���紲4�ӑ�"�vg��|��e���L���Svb�߆W���WP��oT+��0rj�*kj��!����[�����A0�i��N�Z����;�^[��Gi�N��&雗�~�T�ߧ$�>\cz~l�lזy5_��w���	w��9��.S�x�$4�~E�Qa
�r>��h�4��܅�K�*^b��d�?8��Tֶ����d>���8�&��3�>��2W��vvj�Xp�!>ٌ-�oO���'���a%���10��AW��$ؓ[ �,����%��J7[t���c�YAi��f
+(�*��xr���6&C'�)nw�}^�������k�$��_2$�=�%U�������1�;�1h��˪G�O!fy�-Tn?�c�&�&��c����6��r��)_�hSK�s����Aw�䃣_�xS���x�˵B��k6�3wyRHn�^��p����^�����u�'��5�K3����+��;k:S�;?nV�X�fB�����S��90�Ԓw�@17�t���^�fg�{D�n40'����WVjv�BFh(:#���$�A�:��ظpwC'2cu��̚沉����&q>�`�JAj¤��F
������ �9�	n�$v��g"m��=+ޏm�+s�������+��OE�W�j��0g�WQz,*��b�ϕN��
�ʰI�
w���G����gffĭ�h��^�9%#��)���J�=�f�N��6C��d���?�����E�;̐+�� ���4�8	��3�C8Ҳ;����F|���3[(ޟ\������g������c��^���.����\�=��[�rov���(�����Au)��6�d�Z��N)� 7MCl��� S0%�Ve,���:�Y��sa��3��L���{&��ߌ��{v 1q��ʼ�fܴ�]A��4>ԉB��r������	�	��Α��>�k�6��f�&���^��:���V�_��Yd���h�v��N�~�6�da+�j��.o�����E��+v���k��Si�8�r�К�P#�������r���+�Y�g_���[���Q;ntJ�g�)?�gǵ�Y�.v��c}�C|��ɕ /Z$�Ci��lz@A!c�����{՞ns�r%T1��״��pW36��<�g\IҼ3u���t̃�t�����L]ڰQ2�ݘe!v�\s`k)���(9l�Z6Y��(?ں����iZ�����Z�7�Gd�}�ж���JM{�y�'�D���"��=�\��f�`[k����{��W�Y�<U�D�~�������z6,����n3��� A�[؅<7�+�ܕ��=[�
��<�ʥ���y�*���i�Eȗ�zng���g�#l�pz�2�1:Q�$aX'Κp�k���=±�΢ҍj���U�P�� +?,w�!�ɋZ_�����N�����	�.���n�W����4�����2���>��\����=Wx��FQѹ��hv� �<�6+I�a'U���,��g�sav"���{F\��b?�*��{����[�GY�e��pw�����1���n��N�տj�-jƂ�:���-1�1E�G	�ÁQ���e����ʆ�w/�-��0�q���V���:wa��g�|����y����-̰r���t���`؅FXy�3�����sЧ��[�;��X��Hk\�c��>�<=ۭ-uA�1�I�J�x5�a!U���՛{^�Y�e�3I=�w*��.��i�?λ�Af/QY�7�%3~���yv5I�[W\G�$s����4�~�RWUH��0�
WCZ����G�������̆[Ƨ���	�[i�-n�GxD�n�*��<u�H�5�\�;�\	�{�z�O-6Em��j8��i��ꍍ��7Ű���͐�����E".�Ń�:TdCqdy�����9�2,����'_uǿ�TT�H.����_�+����}��Ӭ��_B�յ��4"Ʋ���"gB],1���x�'����)� ��u���)͹�Dϓ�5Ӭ\]�KO����%�YM[�3�	��)G��:J���p��L:��%�c���Q5"�9w<�R7A����xn٢����"��+Ո���5f���@�8B(b�2���p����6�o4���\���@̪��/���<����f���w&����a+}�h�ڔ�m_r�I��t�%��3hG�d�Z��u�p�˩�2��#��ۻK K�>�qK;�D��&�i#$�E����V߭�'��*��*�"-���h��t�A$�pC>eU����p��Ap*�{)����2W���*q���3ޟF7[?�O	�C]\j��t=��6����ͫ�����X^k*Ə���,��\'c���B��M|��ZJ���`as���'\�nwvb�F��/<e��A:��cU@�2��=/�g�x��~2��8�ֱ:a}J8��g�$��)�����m��,V
��2}�'���b��@=��om}Z��έF��F156�[-'�������}2h\��?١�O�00���g7���!�5����u��b��)�+�$C��c������ȓ�� �ZD�
�#�g����Fr/��u���(T�:����s�p�[����ëa,����E�q�7�$0j�p��H����
�Ȼ��OZ/�v�*W�^��5�[�B���	�6���"z��cR�1��XB������j��l�<�� k�/l|�t#��W�͎�,nV�y*�
4�Xlۢ�$��U�m��}MC����_\Ot��������>��g�`���b����_ʋ�\�ܸ�ǯ?��Hx�Ny?dڞ��Wu�|�Pc%��F��;f��.E��ty'�Ɔ����|D�M:�㔗�_�e����$�I��+���,���̾s�p���e�k�$:|LT�C�K�)��������o��.�| �flՄ�29o7��Il�����s�Ћ�d���zM��R���?k9�'ö͘�$����M�5i����[�����'�?�@}��m�w���K�lbkŹ�w�l.�'�A�W�?�S���>�?�2���0^<���%E:O�뭁'�Q\%�%��j���x"�R{�a��w)��l�.�3=ny_��H��	\�Sz�����7��Ч˳��\���,��Tm��f,���V��M2g�p2[�'�������
�N���Ob�/��C�/����k�3����>xŖ�3���(����e�����6�3{4J�/��h�iDy_��ʈ���W5��9�X���D��7��2_��h��@;�hh�9�*	`E��@�X�|�H֣��+M���1n0��͹�H�|�E(1���v�����n~��D�m��Ʊ�4�;�y�>Kt1N�n����=+��Ý�e%Ohбw�vk�Ѐ7�b�b�(�򂶵RYScH�Ϯ��	Q�p��#�zV|ZVܼ�;Z�`�+*�F�ɩ|�%Xd��;L�����ӵ(�! �vM}X���\��X��yJ�����u8���6-_��x��s���4�D����[��1'����hc��%�ធ���&�3d�sx�1�W̧�) Q~F�V���m�7����ϕ�_�d���_���z3N����v����q�s�-�V���d���g�+jڋ"ĕ���=h%� ��B�A����G��������HG��v�5yq�-7���B��r���9�I����)j�l&����	ξ�P/���C΁�sXP��ŖI��E��9��2�%'��`v7H_V�{ǅ�w�L�*�Ɣ�>�t�<K��g�uq��*nr8"}�~�{+\es12��T�I�8�����8���qI�Ut��#+�5�y�wv��k��0�O.�n���V��l�//.e�r�������r�$�Ɨ{�!��h��.{�G���r��?�]ޣ��9[�Ns�[�_����);�:,��j�4��T��~twy��ΐ?�a�r�t|t*��{<ud ���t���]�n����E Ua�_1	�C)ف�b��]�Y���n��XMw{��å��\��J�~����$S��eEf���9�S�ɗ�M���/�>�I^)#gI���=)p�]DRyV���sW�ĩ�q�IasZ���u.�Z��a��X���Ј���c|�b�O��K7*性��e�Ҿ,k�0䚥�|A�Ҙˍ�}�KU�t��m���C�KЭ)I�'�5W�}�s���9 ���=���[!`�7fA	����*�`l2��T-~<F�_Fh0���%#)�Ά�Å16v��w�������D�Ify�C~�1�JxR��I$T��	���<3zv�G��������ox,��{pPna����5p�υ���ur���AXK^ل4V8@��79�B�X�&^���_PV�ۥ�9;��&�Kc�'������S��Y��\����jc�*I0+3V��g�j��K�g��]8!B�E�	p�7�m��<Ί~zlɾ�5-�d	����O�YvM�>�f����靆�Ew��[ޭvܲ�-WbouZޕ�q���%� nWҬѽWW�������,I��w�Kw 9��=��[��2'�xbdϑ�������* ��� ����������U�c��IeKO�|BN <�4���q����L\��T����2�~����^8�q�.RV[�<���]`!E=� �N�_�$�[���,������	<���ht/`'���e������R[�1�-��o�"*�N�k��+���ٓp�D��M��ɕ�#�g����vY�VW�D�����Y���M�B�$��W����>w�a�(���T/@`���B�84gزeTΑ�K-��.ǃ=
��c�pT���vt\1���5�g]�������G\�� �}7(7���̅	�n���"�9��/��ik�/&!`Ӻ,���,v�����8ƍ�q�>C�'��Z��P�����J	�zG�?ˁ"�Ν�#��9-�-��R+�a.G�}3��2u8��9�b�_	[�p�8�H��-�[�C^���nX3+��9Q�O�o1G=w�J��[�F i����~���PB����8��F5�V~�:�b�t��Y���e��*+������Љ�Y���=^����`V�O	��+��X���
+�]$l�d�������� �� ���Ȝw;�pI�u�7U7�Hw��{�?�Q�ʬ[���/ex�����q�� W�vؽ��&<z�o���ۚv�[=�K]�]�@���Eӽ�_^�<��>T<w\b�@6HÍ/�I�V�F���KGW��6~�����hi�*	\��u���uM���Ž�;��4_�Km�XMz|�)[�[nN{���O���i+�/z^"a��~d��L���#ٺ�iC�}o�<�-�W�N��;8�}U�ÅS�����7�3(1�z#� -�����p$W��.�����H�AK��Mn�`��bO�4�1��ٿ�5������d������p�4s���Ɖ5��c��X{�Fi�cc{�:�B�{�fc���[ �p�,ꅘ�G��L�W��	~k7��|ςڿ�5~��~i��D��������Q��2q���mA�Y�Wl���ӳ]}���(�)���z���_W�p�IbJ���U���U�}q�U0/�n �K��O�/�e������zl6�n`	N �iE�03�@r.�Pd�+�b��í������e�5}�ajby��z��!�t|u�	0�+\�ѧ�~u��eV��i�3��ox��(=��V�o��Vצv�f�㯱Ʊ1���6qS���k�h�� �+\nmq�r3���/�d`������[���ڱ���B$���~��k�Bx��
Z��źZu�W3�r���σ�m?��Pj�=[;۝nv]{>[e����f;I��V��4b2g�U�`M���&�ľ[Dk�����d$�M-������A �\�����ѷe��证j$���^��gU�&� !�&���Dk�@��}D��ٞ�UبF��!�Ƨ����m��	�sL[��H��I��W��Y�����*EA�X*5�a��{��u�;aϋ3�|ˮ�&|��r��HD
�k�fp1M����4�,W泛��&)�Z��;nEn�,�­����	̺�I�6&S��	�gA�D+5������rL�mv��5�|Y�_{\��A�s���^�gG��h��}P�]�W8���Ջ�5�*��-��'���.��Z���s �S����Stt7�;A$#��&�u�G���[��}HT���(�!L�e/Z����H�_��{���%ԇ5N���W�IyI��)Z���O��J�b��>��������R�K������\Hn���z���G�}E�ihf	��	ש��="�p�Bu��B��]�pX]�y8v�/�A�@����X'�M^:Z�r��*f�T5�@f4��!�y����d(�LĢ`��a�k��b�+��%�+Q\DfT�e>.{?͂�
0ک��J���x����8�ؚ��3*cć[c��?�A*)�����a�������6���y�A����zE<i��U70!��I���!4�Hw��4��ݣ�;���;AGN�ֶ��M�ogg���X%955����g�(�x���0��q��冱8X�z��f��{r�>_��Ķ�1��y�m�`a�9��lH�8D[ϓ/mh{>�$�����ً���Lq^��ǒ�t��:��.�3�d�Ę?�K�YU����ԄҮ��'K�'�����-�5�D�}
�t�pC�'M�0@�"ڟ�U@\$~EĬυ��&W�b�����Zwor�_����a.{,�z���zmXJ��,��x�˂��cr{,�()��I����}��'���[
r�OCK?Re�~���w�N��-s�X�&�8z�h�~Gơt}x?�v�wYg=�z�u�"2���%;}D��l���~2[Re�`߷�RjWjk�8�FiP�+N��5i8P���]]t<%��z�&�3�P�]�4����׋=H�֘�hW�E�c�p�/��ċ��˼��%�+;��Rlۢ��CD6�T4�2XE��o����t'��bg�h�Xl����<��J:���o�S�CI�όJ�+=V�.���Bw�b�I,O�gr���,끫ID`۟��@)�걟͹��1�[��k�u�ہq��|u��|���A�A��W�L��T<��ٟY$�B�7�ᔔwDVzuYxqx�A���dalln ���d	�'����^�-j���޺ݤL��{Pb@n\��6�Q��+e*TI�Ӓ�H/�_)����Z��p�O�����?����܈�V���b7ĵtcW�Y��6�9�Oh�2=h�u�F�a,���I�K�cZ�c5����s�I����XD�5�bHٟK���	Q�b��PA�%lXY�tg��c�S~}� ES ���#Wd	S�if�ķ����gY��I��\�
}2S�R,������P"���F�(3����m=���"���ʋ����Vg�~�{�����j��ô��?����h�"%�������Ę#TqK3�K�C��B���q�so����p����v��,��Ĭ����?+hBK����>�Y(=V��MB0��g[��r�Z�P���8�L{��|�+�'��;�98���ߣ]�3 :,��7����2��*�ڍT�	F$.J��mJ5���gJ��zpaU�zs՜��\� w��M�֥���Y���kL%]Ms�?{/t�7�Z4�K%)/��,!��|B��~�y��p�)�F+%�6z�r$��y�X�ȫ�osd��"�l���7f�V+N<&����q�q>!������*��8���1-`Kx��y�&�{�)|�g�J��-Ye�[Q�L��;K��.=�����G��$�3������
�hV��n��-������+ss��-m�o�a4����v&F<ݘ��vۍ�ia{�U)��g�	,�>D��f�
e��gPdVSp6��_���K�� �����Jf���7��� ��6N:�Pe{j�
�/�B�>��p���~�KZw4''��R%����\)�W4'~���Z�.�}���E@�_����a�=��A�k�>c[�4-n��S�؋X���{�x���a��4��"�7g8
�L��ؐ M��B[��VB��#�^��b�5�s7\�U�c��B5gDh�\2l�V��<�U�p��7��� _����*����-�m�Fs31R��5?�:`_��.Г6!#�@������u��P��xNω��$�ʸ(�E
��г���eɓ!C�"q��z�V��q���A�F�����	����?��ݒZrx3fV�s� ����5R y�@�������x,�&����Q����	5���#�~�9Ot��2��_��ܘ&��_�YG���"}�'�k������_� ���19oOv��YX4/�98
�B��g���b5fϾ���:~��9r �qB����'1�]H��b�����XLL.�9.Ķ��g:z�����L��R�}������7��4~�h�Qi���[:+�#;l
�|��q�������2}���W�c*�~Fd��5X����N�#�B,��W���~��/�����P�.��<׊�a��;XeM��6��� ���XlW0 Ӫ6��U :5����gV#h4G�!R���lc$`aʾ ���ί�u?���K%Y'$���>S �	נ䳺`ᣞڎ�`-�w;�A��v ����F@H��f?='��׆�^�sꏕF ��p�e��N��]����lWИ6Yʤ��
�@<*��ῐ���޵O:�~WR!i�1Uv��WG������ŉ�z$�n����Bj����o����!����ڔ?\�ߴ�] c�2��O�P_䌏{����ϟ]��0���W�7�����I���څ*����!�!c]���7zhl�j���	��R�A*��~m���^*�a�+��>�ja(���X��NX>�N�xb��aA�`t�.bsz�:�"����^{��;vZM_1�Ç�$�vL�� )!�yc5}��W:��c�JM�k�����VV���27�t��,[I l�sr���q3�Ek�f\���Y�?�@"�2�T$�Hbig��=���.�L9�}@-LLe�DZ��^�#��O������Ո�w��v��2� �~�:B�-3�^���!�ԕ-���`3��C�N��"tAg�A�EVY�B��ҝy2~���\�K��㱗,�0{�}���iʻ���;���2b1���G�ҿ�ʹ�8�?H�r�GM��g���	�lP�  ��/�/z��2e�^��3�$gj�K�8-�N��2.����ђ�! �(��y��&ǞN�{��7�ק>���ݍњ��[�æ]|�_�tA�����A#]Ɛ[*w=,:^~H�G�A�gr����a*�űG�mZ�g~\��^��\�H,��4~e�w���rqȺ�Ե�ޱ��R�F�`��ɦ��-`�㭅����3�t��|��}B-t���G�I7p��
Vm9V��iaI��?� ͋���g��_5�����cn�1u?�����ňk��E���q���;@�e<S�_��O�Hh�U�ڔy:m�@/V�ߖ]�O����RD탣n$�J�Ԉ�u�J�YW	���=��6��Q��̈���e���\��=P��[c19���*��z҂� �:�m�ҧ�v, ���*�2�q]@:�va�F�K
��E|V��~-��F��i�ࡪ�x0R��ߊD�Ws�`�F�'T��|���������9�r��_�T�~����q,Q,r9G�����w��I>�G6���K�wGD2X].��ĳY����Xۜ���f�z��K��������!(?|S��x����oTR�"��~�,�߆�Y�{_�l��07��CQ֜�ќ3v[n8⫆d)W��1�m~n��;�������X�]@��8���m�{���x
!�|Z7zHsQe����o�14勃T�����F+Xح�v��>����Ԥ�"���c�i\�-�����y���ZIM�
�������_�UEG��	���Dڥc����3W��F Q�)nS�G�/���e"��m�tj�c`ﾮ-�~��%1�m
��o���r25�'y��9�~�S��\�$�KE� Rlc|��{S�Ŏ1�lًjĤ��X�ъ���N���1�]J8C����G)�=����ym���Q�0+��lϧ�+����9�Ɂ"Z=Y��8QpLR%����p����6�|��s��Y�������kr��L�Lrr+G߰��߽CB�2�W�/����_?����o����^�I0L)Zcuw�X|�?U����x�0j!-ꤐ��BOc����\~8��h)����~�_��&h;�b2�F^">�^&�,3XW�����,�+ݳ���ʺJ)�'����e�{z����C����P���t/K���Q��������~�:��
U寪��^E��c��4�l�P�;Xgs�����ְ�\�&?/�t��I`�t;>f���s4�cz3Br%wЬ������QV2c�$T�$�����NםCKM��x��ȫ�Mޫn����Rm���n�<�:X�@���/�L���r���Dkd\�hT�FB�p����"s�6 Z����}3Y��R��j�<Qـ�������ρxڨy�W�C�>+�E(l�\-��"�D"��k�Ir/�+E��}�	"3��M_�7P�ݔ1�	��	&Cz�߾$P��^�62z���xȵ��/D ͧo�d}�d�4�uyV>z&v�%3��:!��t�l͔ä���Td�sR)G�l[W���bF]:��O���Ў�L� 0Q��2�6ti���D �q�ُ.�������(�����Ŷ�XZ�L��aX�z�|AV㩲�4w�q�@��ƭ�l��¥}'��~��i���D'���A֟�i>��l��<��U��[��cK� �,�1؉;O��r���+�����0!�lOƇ���F�R���d�k�T?���jIEK���OC�a8�H�
6S���]�b(x[-Hx���Zl9�������D��t����-����ZjQ5͏�U�zjuOUr\i��1�H����U��/	��	u��ʿ��݅#��f{�J��dY����J ~qËuFT�.f4#K����C<t|,�� ������7� �h|��7|�q5>��%~��IX��j��e3��6#��0��+�2�`)��i���l��i���GL�Z��cV7�~.�!k\�B�X�4�����S�4����
D]�"Zfm������zڲ�4s?��L��9R*��=\+�{o�͍��NԈp���Á����4�rk:@�/�m�1+�8@Z�J���%:]��m��u%ݹ:�f�J���P,�g��w�����?��/8��
$��/�ВC*s�vI}ޯr��m)���J��w�a�e}.��=�?���(ܗL�4�� VZ���y�+oLH �76� y�jqzv6�?�e�y���"��ӂ4��ܭ��uɛeR�����ʅ�c�}T#{پ���'� Ӟ���H�)�T�}��B8��)�e�B�5�v��/�U48ca�6�ue����l��_N����F�n9d�t�K \�-8�:��lܤ��!c�G���p#�Un9���&�A
����j=�������� ���9�F�$����g�б)�}�]���(��7�m�^�p3ت����:�Q����3��Ǭ�r	8̒�J��dpfSV�ҲJv����/f�3^Y�rq2� 9�)��εÁj��ͨF�X�D�xg�x�^Ѣ!*5P���&��f�8A��JSȟc���h��y�*v~E+y�o�Nz�����z����QVg*�7��]�Ku��
��	giii�k��iv��7_"d�9Kq�+��Q<Ԟ�}]
Y'm`�S�X�llLj?&��lq!�%ߡv�F�ū��7�6����66��p�z�Wd�⺸�_�c�2F�61���C�����\��ѯ1pCg���q��]Lx�b�׊��y�RDR/qa��NI��]H# PV^k�7���Bb��,���t�����2Q�|}��Q�����5&���$j��R��4�x�h���.�^�"ۙ����DJ�?K��&>������7�,ٓ�h\Q9��"��b�&�i���|���)��<*esL?b��t�����M��t7�س�D]R"%^$�����u$[泐1w9���YcJJJZ��X�.��n���C�S*
J���᫩��I�u�U�����Wڢ;�����DX/�Fk�rat��n�g�z/��{�~�t�*>��NFf�"�.�����B�\�jZ�1l�#냳oT�_t��ĥ��j?� �vM^_���`�u�	E�H��n���u�i�=���X�0��E��9k�}���i�h�*?�3�#������s�L��x�N��U�<�>C(��U�eV�e3X�[a��O�b�Ⱥ��l��}h�q���l�����D��W�S
T���GվsS��]��+Qn��/�<�p�5�Y=�g
E��sM� ���vm�h0�)Zs�t\N��5�@��K_���kV��_�w{����X�}ץc���7V��cV�b7��2?���,����Wc(��*6�j��^5���C���6`�[����=`� |�	��z�D�}c�6�����ٖTLt�����]��<��Cm�Ƚ��ݟ�,��RL��b�doTc�C�i� J����b�(G(_-�p)���͑t#A�ߓ�W���s�Ϲ5�6�޺�E�����dm|{��E�U�.+��&4�3�\ �f�	����Ⱥ"O�P�%�:D��,u_����E��e�|��2Y�
]G)�7#�H�+�>k�= B�-�����gU��շ�BFm��kױ!`af�wsy�����9�poL(��K2��lݪ�c��M� I���؛Sꥇ���$��
�}��q��움]�b5�,Vd��O��)||%###^$w��;*v��cT=�(�4>P��hP�P�m[��h��Jv�>g����[��tq�Zi&���c�W-�iR���
�$ҽÖ��]�b�
�
�,������5(>OMAD��-�ck��qt�Z<��f��������.��O��By��8�A"�6�:)�?��w�>���wz��z�O������~"�d�J�u.��������'թ�n��谏`�qJw3���_�A��I�>�~�mBCH�ɽYEP�,Tr���]ѐI��>��7�ma��%�����<�d�z�_!lT��Sseh��͒��,l�h66>q�$V�f[�� o�nGm/qQ������]�tw�����
?�V�<��� ɕ����@/c^�q������P��t���z�k6W��9�?�oovC�CGϐ�Y�7�(�z�hL�W�h��&qy���=����=����>�6�,��_?Md���#Z!�S!����5�Nf˟�G��q�Ad�x�
>|�>���@/��o��/v��6��I��^��m�-��ԈVm�	q;Sn�o�e���K���d���4�X�~��#���)���]��#� �ˎ�8�Rko�9�W	�b���i�\cΓ����KY��~�N�D���c3��H���41k��y��P��NZ�r���!��m&×N�2��J����Dm����B�m)1�o/����3�^[��Ϩ�?$��?w��m̕@j��΂s�f��{k�U��n�M��y٪��X^�F,��'̸�0E�AW�~[�˱�LdM}�����5b�O6z �AJ7�V<nVS��5���K���������n���w��M~�|�o�˳&u������ժFX�@v*� �|δ2��Pwl@��X��y}�j�(�_F����+�$�
)���P��E���� �)د	^f��(d�zp���a"sJZ�;H@������%q� ^��~T�̴k��)�t+�uI��5A����smΨx=�Rl�(D�� :�1jU䡴��0I�
ko���Zu�<"�L%?xV9�z���7��B;�܋�P'I��جZ�����UZC�uEͨr�����Χ6���mkc���^A���c���6�sRo�=��mE^�HT�4\���͠@�G�?�ޢ���oV3p�����L�&dKK��aI��P��R���Y\d�Y+�W��D��LF��hy�`� {W����wq��1�%@sp`��黛�2��[��UwSpu2�s��.��/�9�,)yy��S�m���W���/��.�SZ)%��~P,�[G����d�5���!�ߍ����?�V+�_^�i'��y��Y�6��?�ߥJ �+�� �3�Yorp�!Ⴢb`��4纾�e�*/%K�kҏվ���ZӽY���O"�"o�F�9��B
�;��_Wԛ-�)�?���$RZ�.�n�4򷌌�,'w��B�E�/���/�B8��bͨO��H����$���(#>oln��Xw7�2�A�{�){�����5�2���gCnN��K������ ��� �3��h�u�*�Bdy̟�1�&����8[2"���`�稦����|b�f�²�ⶤj��i��j�ÙN��_:<f)��|PPЁ��L?i�׻�w�Dg(��fި�Y�?xT&��*x����fi��2�^?�
u�����0�_A�F]�q8��#E(lg)�����v��Ry��M�g���Ǔ��c���H���UPQ�B�u��0��ݎ ������dV)��;eQ^�S)|�g���[&Fk��u��us�ß��8O��b��D�]޽sx���o�Ҙ���j���2��/�-�ٿ����s$<�H����i�!����Ki�\ 
��}i�Ł%�@���Ë$�ۯ�����O7��L��*zw�O����ס��'q4D���$1ā����S�uj��s9F���Q?�g����+��}=Z�[MA*��WN$��0�Bm8�ex��P���W��ۖ^.0����<���X��g�Մ{SƆ�n�Z)�=a�c���Y������R���lh۠�:���[�ڃ�C*�i�!a�Fłr]�A%���R��oVX��x��/�>Y#/��~0�4�H_C���7�:����ٝ�$d!��..ˑ؛䁥��=<{��]��׫a��-�����>�o6s�5ro㬟�G��T�R���*K��G
J�h�;1Đ������"l���9�V������F�B�� Z-vG^������yI���7�GZ�Mx�7;���q
��I�+�`�P,L��J�4f(�?���b&���;.3���Ѯ��W��@φ����pg'�!}��m��ߍf`ApЕR\[X���mӝ���̈́_�n��@*���j�T��DK�!wk[�3:`���Jʮe�N${�p{dmg�q!�q��m�șo�!0J(�vx)3���4������[��l
.顨6���.1!�7I�V��R��8�9�_��M_jjͷ��?��3����{oѓH-z���#A���E�DD���^G�ޢ������{}g�������>g���>{��hM}�nY�0酜�� ��Q��������eK����6��G���	���K
���Q��#���Ir�'�7��?+��`C��c*�}���ԟxz� v4g�KE�&���k��q���UW��q�{���_�ld���w�%2�p�S�>��{X�xA:Mڛ���2V\�]�ꖕ�{0	<1y��o�yz������	Q���6F��r}����u�8Ib���b��م�����9�Y��0_>�鿪��*h}��lh��
v՝���{�a�حƃ�J��8lsL� �A�W�H�8�LM(�F���$�����J�`MQhN*�����ɉkso��RS_/��9ѹ+w���5�����K񼽪�C���_��_��[�P�e'�e�餳�f�����LD{�\o������Ǉ����V3��Z�H�o�>��ײQ!ڶA)<` �ŏ��ɶ��e.�����ן���D���IvK֋��p�ɑ�x)A�/�Zin���m�'ci2����S<��ñ���z��MS>�#q���#ҝEz�p��[���y�r�`�"/dL�8�N���,����n/�t�ղc�/K��zP�����o%��:��x�j�%؍� �V�̠a"��;��K]T7�Aᦱ�;b������P������dY'-L�w�@[:&�����&%��+�V�fZ�'�?�J�z��ٳrM��[���){�Lju|/����K�3\���Nd����R��|�1
��a"�z׀�J ��Ճs"K`m�2���G}���_�䴡ɔX7�*����������������h\����qR �)�/�p�|;r�o��tص�e�ӱɃ����֛�}S���JFi����w�����<?M���-�X�H&]�b棉�.��͐�>���Z.�)�VU�z�N����$�MA��bykC�!���@xN!��E���f�9���4�҂z�rJK����1������;H�e|��&�/�E�ȏ��:��ೳO�<i��ߨ����ӣ<::z]C�C�TPP�<ۥ/.)Y�9;;yw{u�,�E�,���J���#x9R�UY�R�&A�����&<{Ϧ��~G�4�:��J(��ۡi]����0�_Z������|�_��;W�6-���x,�8�8�T����w١׫m915�o2��5o(��F!'%�˼4�A��9�h�q�3^��)횭pt�턲�ؘ�D�����ls��QNlu���!��$D ��k������ ���6ʒ...����[��=N--�Q*3y�� ^���Da!���(ZR�y~͉z�?\@(~���^�fg'��{/TBb�	+�B�*Vf�p?4�ef`�w� ����n�g�ms��g=J�sx|�GDJ����ʿ�ޚ��-���8���%3[�ɯ종�����{$%$F����y���x����y�I��B5�_y/�F����`pBb������~O��^�/t��+�u�10D��奲��i�����^	�9�3$����hu8XW��S��j��X_s6E󇗻w�F�G���kdX���"'N&7�(�׸�n#�$>s�� ,;���|;@c
'٢����`s8s-��gr�3���^N�Bܾ���~L����k�:Ȼ�k�:C�*�Tɩ�6M�}�<ݍ�	�9����11�h���6�|��SMъ3.RM,�$,8rd�F]��6:@`q�b�����n)�*�8�6<�+Y�7u�7u��я�U���g}䎈�.Dsd�O7e��/ ��3����4��mz�m����߸�^������{ ��Zh�|K�u(ޗ˔�J�� E�$)�(��ǵ�Pg���ǿ4�����n��NHBW�=,��k�����Q��T~g����r5Vr#uKR��3?"N�ʶ+j�氧ɨ1*!>���x*>U��jgdW�}�����J�r}�,ٚaV#"j�{Je>{~<;1�jA��H�b.�<Uf�Fn`b�(���\);��2���6��K^K+�y�De4ۏ;V�|���8���9F�4���ϣ�	ƧD�>�*}��S+]3����~mu���ĕP��\�����󾤤���­NmzBB*���F�b�݁�ZZZ��E�s���?�v�B�b����7����yF�B��T����D�M^�	t)
�t�E�.
˰��+"nϾb�2����`�7��K�;S�!X�}����0\���u�{aZg�{tɸi���]�x�}c�wXi�����@c��ø�'C��*󋺃/ͺ�����5x{�	`�H�<id���7�pm���KeTB6
�#֡�6��;l�b���[��H�Jy����&��.���š��''W���> ��k���#~�q.�=̬�U�Q���[m�9��=��'~Y���[��k��D��*�^д�qՊ����e��
Z�3xun�2]i��������S�X��|�w�_��o	��a\�DX�X�%$�n��M�*M��.�ɷ��V���ř�ô.L"�F�	i����x�Z�1���V�m��떇�~r�
O�-I��!&��w�^��={g��=�������#��f���QVW~iB[�;����V-�kg�:靿UL%���AV<�P�_����rs[�a��G)�~����V ��mp�Lq
��ފ��v����N�w��K�t����U.���u~�wH����dSq����,5[=W�hM	�[�������mO � �Q_R�_�@�gs�w]��ԃf#�sw����J������f/15<�?�.&�uc}y�.�� ��NqI~��0�P�c����ٞ��2�S�G� h�AD̊�N�;`������mvC�$������g�˔����|L���D8w������;��b�diGH�N����*�\��K,ܴo:H�ј�^;3���6h��K�g
�C?��u�֨`cUz�jH/��W�oV��+q�A��*�s�tp�TQL#j2�D���̺VfD�B��k�<������W
 ~W�����.1I�T|���F<z�yMb���	�y~ն�C'��뫊�����s/���S����IB�]0�;[8q<��q�FGE��-� �ڽ��
�HL3酩aS]�Y�WߟvA~�6[QZ0�-EO�ƍ��s�c�T�"����s�uT�����)<��'BXm��6����f83.�	�Em`�j�h6�3�c�˭�����_F��/�z���vgy#�	˳ù�_�{�B��/����Y.ꤟe=�	28�=��貓��`�T� ��~��&JT˨`3H�}u�;��η��Q�E��@�zv>�4

S�NK~��Ws`�b���1��ҹ;(���#г�8�$�|�e�0y����&�*�|�'��G4�q��:�Vi=����I.7���/�qŶ	ևZib&����OV<A<w��)t��Y��[_���FD���yH8x}�4BDR�S";P�"n��;���G��X�!��(�:�3͕�(��o���&O'4`O� �;�^s8����uv$l�:�Ď��D�gy�v�����"رԅ�Y�W�i�`���1�����B��|�͟��|��FU�kjz'�^c]T����w�\���?�:�||����k\e
��}�(����T��뇽c�7V�վxϣUU�m�L�x���`Lpv���U_q 7�6b��W�����_<��	)��[�u�����п�-�������{1O��A^�����O�Ž=u��#��?��Q�Q��R�x&ɄZ:��+�Lsh��L�\Z�'��7���Ik|�U���)ڣ�ذ���f��$�^��i21g��Z'�#��������׀���>W�s�7km�A��ѡ�8R�O�D�o7�bv>bk&=A�|I��"�<�m �u&0�랡�o��nu����:�f�KZ��xEX���{��
Q��a�m����C�-�t;�e=EV��B��/Q�ᔐ��8^��g��Sşp^�މ��t�����R�bO�t�ssv��!	{�Z'Y����06jc�q;��.��Aeo����w�d��k���.�:�[�Cm�3�Q	}����-m2ch�n��߶��%�\��?F&~��L>|\�����f��[����3�+"�����(Z��_��Ŏ�	�=M1b�\�/^�(�u����R�2�YvnK�|+�g�T��n�B$��x��H&g����h% h`��D��ﶷNN,�"���`?-��N�b���y-�t�.,��s��}��H`�%����&��ٮ�3��?e�_��͒B< �}7�����; �g&qN	�b�G0��=m	��Y�������q֨�~ei�7bIE9k���'k�F�������P➳���Ew��HD��j&Kxx� ��2ݚ�8�/{��5#A�߰�y+]���y���I��3�}��/�l��F�� �$D�O~���W���J��%�&�?H��Ox���I7��,��+NɿJ� �#Kd�����D�����*j����d��rE��A��	�Z/�}��H0Z#P��3,>��7��DK����_r��,���9�d�L�p��X]_�J�i�ãP<�q\��s�~��S�m)\��Yij:�}rIPyDр�f�����S����{�2�S�$�NZ�Qڡg@@�"/�Ct]�d��t�V5�Gڜ)�i��Հ� Zw��n�z�����q*=3.P-��\���`��W=���,o}�`�6���������"*�_s'�t�2"�y:4�b6r�ik��Ͱ��S!�Ѐ��	�ah屵���Q�cQ���4���]G���!��	�\�%�Q���p�O�J��?/�'�-S�vuay9�*��6<҇�n���!	�d�������9w�&�wJO|Y�$�bw�a�(�y��H-�����|bp7s����@����*X���R{������Y~y6>zĚ Vǳ����F������Y�ɿ� =�(���Qg\�m��Q!+�xDb5v���x��^ ��J��&���j �jqK�fSƿ��yC3(�؁8�Jz6�̕et�_s;���"�7!�uT��C�!6�~�{1��j�H1�����[��;`탬7t?~�>�z8�aq�{u�7� �o�����Õ�f!T�Q��_�R$�<�*�u�z�W����/�N���)��z������Y��&���M��X��3�P�">��0e]�+���00�����M������6/ND�����B%��h��I�d��`��µw�C����s9��X5�B�Z����~7���?����6.`����_��"�1���n�6~�����\�Ĩ�&$�?�U�M����Nj��CAf)�%��r�z{��0��%��ׄt�2���I3.,,EJe56�P��At-��F��4�&gg<����Ʒ���²�EΧ�I��<� �(h�	��$k�sB�)�=$~#���0���7�9�/�q,+�c9��ʹ�U�.��/��E�S��0�P4wa���n��mFU�m�b�>9n�ց���ި�@a�����(�P�X�l9��JQ�B�2WJ&�������L�H�>�ϐ��]F-�9�{�ɾVR�?:>�w���s� ���r!�|:�aS����d��s�rR���S��I�Q_�L�yc�)M��i��n�6f#iqȘ��ܙ�bO_���2�����ȟy�8��V������s��fۤ^�|��Q_����*3�
۳��8���6#�Gl�Q��t�����ŧʋ�:�:�@\(��RS_�s�%+S0�+Z�B-�Z-�d�b���\#eggg%�o�[O�ߖ��&�LG��$A�G����P䯞mb���23GJ�*K�ﶟ2�l7���	qq7r�Q�[��mMz�~ �?�J���W[�"�X1rL��6%㰔V�n�����c3�=!V�����t�(��.�T�P����uض,�D��6�a,H2� �������vG7t�ƒ�M���ݙ���ȨH�5�v	ʝ0���zT7D�a�K��L�SpGQ>�D�eJ������ ��(�p��1e�9�>��b�N�N�z�N������I!�3c�/zb�<������V��VPٞ2�������b�����5�k����@d_<���N��^GlƿvHRB���#E�Nr��:E	�$�ϟsw�iDO�kp�A�L��±�'W敮����֘�=��;���jHNN-�d���D.�j<e`B�8��ۡ<g����>�/���V�a�q�
��}����FF��O���A�^T��{��Xg�'��#Z�}+��|E�m7�ݧVkE(�YG�2S���'7�SC�.S��j%��^�u�[��<��;MJ��A��rr["�Q�u&	 ��G�;��|�;'���s��Ѥ�E��D�����Y��؏�w��O��o����g�G�֢m�D����W(x=���o�e�JӊǙ�������A+}_s�4G�ʁ��D��OH�JɋBŐ����M�x3{��*��}ʇ�b]36�Y�D�C稼OTm�-\]u�
9J1ҞK�����=��l�����ޟk��O��G�}b21�#d��Ɵ�R����KO�o
������Q�m-�����M9/��l�|:P��ނ��݃?<��q�VB�RPT|��>���~۟u <�"����ayE�n��2�G�~�7U�^b��p�s����xr�E�sw8	�����?��ԉ���_F1�����T^ؙNT����^���:�j�p�l*A��o���;pK��("�ݍ�w��i?x3��F4brfU���0�1�ƈ�o�ؒ�� �*Ҭ�b*��Rp�03{�k0={z���%WA󆳺��톂��L�����Ǭ�h�i�Cj�H�M�fǩ��$�t�l�lϐ��ypu�=��d$�ӱ������5�x��Z�4���8���4���AZ��dlޯ�%���Վ%{��&R?��U��o���x�B�)�@(8~T��
����'+}�P��� �AVzZ(�,���_�A!Yx*A��]��d%̹SvOP�[��A�x��k�O�)���@�pLL���LS�u���W�6��im���������G��C &��9���YE}/]�o.$BAj4E�y�Q	�6�2U7-�a�sk�2R��P��fIYV���EW ����wzQЛ�����6����i�䯏��&�D��֩'d��
ˣ�F�P�#W�Zɦ���'Ϗ��y��rG�@0^"RR�XN]ug;����-�.:E��'x6��Bg���{P	����V�y���=���]�k�~�i���Aibrk'��1:n&ߧ��YS�):ByYg�҇�?[=l�A��"�5���!0k
�{�����o��H�[qiq������ɷɩBڃ!������.�.���R�u�X���
�:�f�ĢQl
�� ��Q:��\��[	H�Z�����}	��趤|�P<!�/R+$G�czT�j�>JIύ�B����@�dI�.�ܦ�&���xkC1rw߽]-���]�4Aġ܊��|Yv�0����y֩NX��b*�`��<�x��	��>~�ɧB����$,*�r�܉����ú��ۗ8��O�ASL��s����Z}1k�F���t�ǿw�~KD��t���,nU�[-�c�Iԕ���G�|w7��I�+J���i#�&��5JH�5s��?4���nJQt��uqq����9�T��Nf��C��Ӳ?r/D>�V-�E�Ț%��d�N�3�C�� A��~��yFp�A��9��>f�,kEC.^xA����S�ݩ�&�0�i{�r\�x���ZX���) ��Y�!<�1=	A�s������^)f��u�Y2�K�p��Z�bl�������gB-�sr����!Q{Я^��ޫ?�P�L�'�[;�v��1>P�ѣl��л��Q�αv`���&���7؉���˱�{¶L=�r���zG�ϟ??�?W78��7�<�$����	�gY�\�qss�]ិW�Z��C�E앒��������F�ɣ/����,أ�G��t�Q� ��9i
V���\����C1��A^�k�$s�	QN���,n�Aq"ߖOEc� �k�1w'�@�
ӓ��d� �x�A<��mu=Z��ˈ�A�����:uvO��B��hZ?�:ԝ����m�Bg��;�}̄ǒ�Y{p�S�W6��:���N����4�ߢ>[���QbX�45�KXOZr;M���.U(.VT��K.�z�/t�0�`�@mO$����i�P]Z%��YM����6vQ�te�[e��)!�j+��O��gE��uII��]�/f�=]���9%!&�@9�Z�\͉>��*J!J�za����m(]�r���2B(yG?��c���6V^H��GBˤ(��yp����J���h�/��K�
Ry�!�5�Pv�tb>�R�O�YP��+�qm�,�!��Q�ns��/��I�:��K�n����;�O��~��7�̞m�B,A��"�}GPIU����8�@x^�o!�M�2���2r&&���('���Ŷ��R��'$t2��n����Q�8�i5��B9�)�i��@��(���+7���h�y\JHNOO�@�iT���9�`�\�\�/jӡo("��~�����k��2�����;�o��^?��8�A1�� �hv���w�vr��L��أr��_Rf)Tfv��"����]aP|������@ ��>���y�6��q�5E����[J��z0����o�z��H�/k�cG�P*�cN�p���ÏF�2{�0���5*����z���x��8!�O����xpᅻ&���3...J ϲ���>O�16xB8F�lO{��;$���o�#f�����ΨSk���.��Oz,R����������n�u�;�y����(3�-,@�bY�؏陙{ �:iF_�
��kQ&�E �X�ޛ�n�3�<�IR��"f�i�^���}�V��_��e�(�ZJ�	}Fʕ(�ѥ]�q���A�Z
���˸��QZ'Պ����7*�����l
. #�CAx���H���}�`W]�G�����O�
���ԝK����ҹ&��� �NO�'^�}��x4Y�n�B�syP����ҌVηF�=�q��ۛ�ڦ8�ߛ����l��_tL�F�L2��_n�����5?��`������4C��E-��y���l�껐u@�zt�r�O�b��F�i���Y� �����F�3-7{Z�����\	f���U��pv�_|,
�y�g�<�B~O���q����uH%x���\�Ȧ���*�ל�ڐ��Lby��U������k >%'o4"onz`�n5[;_�n^�0�L�uyyt�8���ߛ�����=IpR�j�K�(�ʮ������!25��R򍅩���h�>d����1i5R&�ht����7��7l�ZG�'�S���pjg,%h�8ǰ��6+	������ag����V�9;p�Y��Ly��,�����ݓ����,�Y�#�a`d<<ZS��	��P6�nL�e�e}L�>#�Û���p3G~G���Q�*6��+0�2(�D3�i����F�0�<k��<y�,�$� �X�呣�j�#�"���ޫ_j�T���K_�#p/6�ŻM �{n�݁{X#$����?�ﱏ^9:�Ⱥ+��r?��OD�ٟ������=��I��8dؖ�ާ?<7���>K]
�۝���z��7Ω�f�2�\{]��YK�c�� ��i���A¶y>L�ub�%�M�1VQnh��.Щ�DW������R��g&��-���>�z��5K$����qa���FIF�����j�_�<Jc��,�aN/���p���1��E��~O�a\3hO��D*��J�[��t6���>��L��V���p֚��Q���g��lR������X���]�m-����c�j�3���lw&x��nP����I���Ѫ�?�����_�u���k;�(%Y�����sbs�7r8Q���t ��P��B�զ���c<t���PҪ�ož�*,N����)����n��`�A�*���%)���3�)*KVr�E�h��W�\�=bz�h㽥��!HK��3���%��@)
1�u�wWz[E
X�L���8�&Ys#�1%uT���Z�˞��-G�5��|�5+�k�7�=#O�V�5«+_+�Szn����t�$WnG�<��Ep��V��D�;�T������7�3��U��J�C;ִ�/B��{@�����ܢ�vL���0�S���u�^�%}h@i�Tpy�S(
���$������
E�Ũ/��<- SR����f�qK)j/����/�T��Y���+*#�0��C��0e}ߴWs4u�(�s�&��B���Ɗ�єV;s��ot]l��(f�����z_m�-T�3]e���B�B�,�	7j�@��̀3**.����@��`d����� ����2.�Mǰ���>��6(�=�1Y�5!y:;�O>8�P~K������k��Q��@v����T��9���^%�z�-��4xY%��:� ��c<��ᑛ46��!c�;*�V���[��J���7>��ދ�ܿ��2w���h���u��7EGfS�IU�,���	u�t��?[8��<�b�zs���Z��p?~Y�jc#37/s�&ݘK�����ڴ"OZ<���C��q%�6x§s���5���{�
+��qI'�凞TVLD�'"b�nGF���g���\(�1X�Q�p�����,hS(���u�Л�P�*���[Z�hm}�CU@��-�^�Dڮ��ݓȋl��ǘreؤ"@���Y�r�������gi����.�(����}�G03����S��A���)t}�#��\��N}$����qd��5sz\[�����K	���Y�~�dU3b^G�� ���{?^]W�X�3���x����b@�;�k��J��&d@+F��$�#���&�C���� _�@�0u��8"P��ٷ�?���'�*�#`#��L&��	�ΪA6J�9� H�ğX��2���MYږvO$B�Y�'2�.C�;��Q:Uܣ���?pFm�d�h��ɗ��\���X�o�����p�!"��&Xwn�����&˹�Y%�0�`��)G9!X�h��C�[���_L�R�,�Гף��n}S'I��(�D�P�e�M[��]�e��:�5�����`R%D�cgVN�������Y{-pr��<�WC��sd?2�E���H�l�'���w�����c��:��^��fӺ1����y���p-9ߔd���D�z5�7�jQ&//V▩Ǧf��|U��9��Ƚ4`�ӗ�b����[o�S�������M����-s�[,WX����$��1\�!sz?��\�؅�Q�ϟw��"S���[
��u�9f��<g�8	��8r��r�ݖm�D����J�,b��%�+�v�8_Ё�}ű�ߓ���Н��Z�N��h�"*0:���ھ@�!�7�$;�:ǅ�H|c$�����r\����?��A���4N�E�&}nh�V7�>f���Z�̗L��� �C� 
�芧�FȪ�X�����c���'>���~��4~����M�X����#	p�c3õ���w���p%#Ƕ"7M�ьR������͐��x��j�]h}*��a4����l��P�}	�U/[����xS���12}��_�=��d��˧����1[�l.�5^+}�2�Q;�Ȅ��vl����:��׿�w�qϨ�z����ͪ�,�������;���X~K���T�R"l�_�OÓ�o�L���m_��9��b�v\�L�5�ҩ(� A�a���FU�{����\��O�N�=��p4&t�kK��N�%��Z!B��&VP�����tx��"�,��|���ʼ�m]�+��7�:�@�����C���u�oR��PvOZ����+� ��(��F���"U
� 8�)8/w� n��:lZ��	��VwJ�Mu��tY�mf�o���"�:I5]?�p-���H�E��g���eyK;S�w�x�SN�����^9���~���Go��A���b�����>zm����I0Y ���冿�H2%���M*�Ŏ���G����(�lOk���?`��"fu�8\�E��w?��t��c,�}w��A`�&1�&���\�~�G�r/����H�4!f t�4�H˒R��}@&q����ݎ�.�C�<f�ߕ])���(|1�	�1�$���8��2mq�s�}S��5F�J����V �U��m�����?��~oetmm������� �60��I�9'Z`\`����{κ"��{~���[��N�S��[ y����yI��U��!stK�����#)���Y�$��)�(.� ���%��*dF�\���2��'Ŧ��o�޿�0���!H-&��dڋ��Z]���`$J��_8��22�tiL�T|��_�_������ݥ��7�,n�o�Ϣ�� c�� ���ȸ�����'䖎�+Wq�A��}씰��?T�%^V�E���Vi8�w���ʠ${����]� �Tq-k��6{��1Kf(o���jOk�aaM��Hy͛m%���T�7�Ӻ�[pGa�����b�8G���}�o��XX�|�ú�+c�+�Bfy�>��N1��5O�,e<�%��hn��^7]�8z��x�2� [���x���T���oy.�K�|y4������Ϙ�.��]b-W�S� %]�do�g9V�{����N1�����Q2|e��3o������%� �7BXs	s~D�vy`��^���إ�Ҳ�e��ܘ3�{F�>���/��>=Yߜ%y����%=��Z �ƌ�=&����I�ܽ4����[����(��#'N3ÖK��ѣ���r��?�!���O��3�6̘2"�Cep��/�I	x�qvGv&�����K�犜��Z�� A�����^R析��t2�l��]�f�݇W���Y�{z���*�>YA�jΏ�~�V�o�lk5ӸO@�m�&���~k��g��/��f�SU�[aC=�~�o�'����k_��,�0UiҞv�o
�%e{�-b���W�k9E0��l7�9H���E�o��dR7�Z�@��9����w���(�&)�ft��P�����'���Fe�N�<i������1l��*D��MM��W�,�Nx33^d�4 ��[�6l[�l���ħdsqL��w~���f����'Wo��苆Z�N�&��,���$PH��^��ͻ�<���Ր���/#�R�0#����X�G9�ԫW�m�ug�4r0C�y[O��F4����4�9s�%�,����2Vh��I�t�����:�A���[_q�y����Gd:w?yG� >gA�d��v�Cw��! G�	<'U��:J�/Ѓ&)q�Ò�l|Y��mV6��T���~���yt��y������
	E�`└��Sb�FS-��T0g�M`���c�c��&���v�w.��,����b���̴�.�Ż<�_��S�`�?�C��k.A��Ϟ��
��B	��cIᘙ-��.��Zy	¹�f$����}�=��e��[����Ãe��÷UUU�����7���!242J��lq�hn�Ӻ���ly�`�9�?�a����y��筨�����"��b�����90�����J��[�7��������[1������y��@Rn�*��0�(|�z�/�i��LE�&�h_m�O�>:j�h6W�3=3}{Gǃ��Tn\�Sޤ����u����9����u�9|�|qd�|4�Z�!��z�[�=�y�kr�[���]ћT�?ۆ�����;��B���5��JI �d�
�=�7m�C&�!����＼�g>�揿�I$5Rb�/�y�����u���'o�!�n��q�|A�r��	o_�☲`n�880{[�'�o)+#��<��o�_�Ei	G;���n��}_i��q%x������ԃ��_v�x|y���G��K��Y�V$�f|�[��Q�u����v��ʔ�Ge����_�DCK���c��ż$���jlj�éc��H}���Я�׫����{����o=��yX��X(��{]\[]<F�w������SG����F*6�܋��[�~8CC/*QLW��m_aʥx�o�Bg!x����"?�����SR�H�oRgG������K����,�e��/*���;L����F����ˑ%���)K�<*���R�o�>��j��lo�V���Io��IYt�xp%f�ڴ '{#�%�"d��#JE-�5Jv܇\C�8y� ������D$�9y-��|J�����D�OG$E��n.�J���VzY��67mm5��6��SS;GG�&���]��.���1P� ����K%5�P�g���yg��QW'RS_o����R^Z�ty�1��Z�x�)�@��P������.��8A9 ����wB3�xg���A�|ځ �p��W���Ʊr��֮�Q�瞔�5�ߚ&�h9�!�E=P���vg�~_8]~�3�Ǽ23Q�y���n�!�ڧ1���y����$:&&�=C#�{���
�&�6�_G��>&l�M����{�p5=����v�j��z�[�g�&��Q�wr�(���aPe�����b�%܋!�T�KQO�0G�Ƥ�`���^v�Q��;G.C�c�y_��na��3<=g{�������TS=�444j�k"��PY�B�¬�p�����:��{�T9���p�o&-_?
�O��֖�I��k����o��˟��1?-H��1�ܷ�ߍ�2N����l��^��������%$V[DSK�d����|���"έI�9�?��Ӣ�iZ��W�E4�?+��'p3�y�[4�N�����»0J�j*����ɔ�O��{�z�I.T_Gcch�e�Z:7�v 5q�MGs#Ύ��DWـ�_eA5�z�7�f����Wv�%�8�(
�ׂ���t#�v4|}��(?(p���XA�-���>8]��ޜ�����>kY|M��m�<m��#m$���4�{�,^Y�̔��eE�sg��p�ͯ���{�����V#�sI7��7,�S'���Lہ΋��4��_e+/���H��_]�t�9�K�<g?+%|��\����Ua`1<ʯ
p0��9ğ�y�;��ʩO�*tǛ<88辣�8��;X�L4v��z��n��q�~v�K»i�C���$Zv�RS��P{rޏ]Yڿ[_D������'���[H�D��Q���G}���es����=z����676��2�fAߞ~�;�����!11ۼ��{�G������ȑ������:G�h㤠�!C�N6��W�^d|��֎���r{�//�܁555��ՁD��0�
���P��H
G��pi�pm��m�Rs�-��#QQ�bi��0�g������v���}�⠼�L��Y�-)�́��X�:N��ꣾe���*@�Q�'	�t)y:m�Zdü	m;�J)�b��U��g�jȪ��*��)W���-���?ƅ�� #Ejs�gz��j�����6�2��.���|�����G�B�p3�˭7�|��������//-$��`�"�u��|�)�n�,�]ˍ���G�PG�9�,��X;&���|݌�<ވ���2����ν��0L�R�2OW#& �ss���j`oَ��/��e��_:[��.��i%�z����������-��n����{\�ܭx��˸�G�ߪ�5�T���gf�����#c�Zh��z��S��keg׏v�U���]1%����>0W�ӗ�s���`5�j�*9�Ih)��^�[��|RdZG@���	��j��ׇ`���5&g~��^��[��u��X+��6�.D`�j�NlM4��6����H�O��P4�I0�+�a�.)TX�{22E���ھ�8��,sNJoI�,�W�|�w>� o}�X��i�Wo�+|i��H��k��5����!�<?�0��ͧr0 �d�e�06��	w:0@EM5�������|:p<��〮2�09������4 �[��B��P��V�ǝ���@��]�紿��|fKۓ%E���J�|oFH^35P ��=�iqC�H�G����ސ�VJ�;�l
v�8?(	��k^��<���s�,U;���8����S����HZ�?k'I<��檅��~OzoN���
��%I��3h�qO]:|ll�B2��H�����fpa#��w�y���"9)��&�4%+,��x�t�lxU�ҹi�8���	җ#��C��Ȣ���]n`z(��?�mo�	ò�£*�	�P�+!DVU̓�����'a�$�±����"�bn�L���y����_�.�u�e��ޓyΆԅC�_��M)$��h���u^�!.��!0qM���LF�0�� �TS�)�z�sű5�Y�D�{�����F�k'�i�X���_��xć 6��rź/2�#m��쮞�a�!!}ǡ��M��ݪ�-��TH��Z��;�P+؈_���䶋�8Q��#�8QQ��ُ΁?a	b5�_��e	H6.��?u�ם#�Sp:n��u
�yo�ݻ����*8��E)HP������)�-����+�q��"��ri�����M&�ZC}vQһ��e�?�����S�Y�w�O|������?BN�O�Q��¹�$]Jٵ�f�/˥�����9��+s֕g���G�u�C���J([ȦP���EHFF8;��l���PvI%�y�93�Ȏㆽ��-�������p���y������~�^�.0�7��N7�t�TE����8��?�Yp��ޝ����~�IL��'���wg�ݛ/�Th܃邟�"}<��N��Ê_�M�b�H��\��m$Dw&N�>���t!�7Bk��G�]s�zo����DQw��D;tO�+�5$T�A��/�ۏw;���
�{n�k�.���!<b�m�584� �c9�) '�l���
K�����<*�k{<㩙c&X7@[N�8%w�5n���vi0���:�����C���oF��I�S�3=��{�+j�=��OD����t90���qp+m�X~��lA"���:�y��ݙ�!�sF��_*u{8��gu�*]W� aY�7|V�u�"�S7��CL���^�Q�O�>���,�~�'ާ��dgm�3�+�fVV�}.���O�);YӉ'ȿɀ3�;�wr�md	�̷cy$6���(��~oj�&���Ϙ8���|��.)kOK�m]�$KH2�Һ�nv.���i#���%��fb����srU$�i�R3o��~!��7���P�K�y�d��U�:zs���~���/R��v���:�X�A2�B�ٹ 2]">6��ٌ&bd|+W%�Jbbbq�˳ Kl@�T�{
�%ꅆ�Ʒ�P���_��`�*b�[?���(EQ1qm��[���R*�a-�~���<[&3qa�q�9H��m������s���;V �N��fu=��=o��3��%����1�ئh��LȊ�VB�b��I5�:�${(�*�{�ݫ��N$θ�q��+S�@���n�㌑Q�������j�/Z@��|.1,���.����-�y�F�3�H�����������mCE����dM�yܴ��7���Z�]�D<?��M��Z����e�JN�u��>6��(�ǻ��6ҊJ���Uq�g��oS���bb$��Q�]Vv��^OZJ*�7KB^bb8��}�e�3����ܣˑg^���SԤ39{��ki�o�_9B�B��8^>�j3淍2n�{����N��������m�Ý��t ���>�QB����_׆���SWpo^x�d�5fl� �"����#�̞_zd���&�;�Ւ�j@^ �9���ύ׀Y���"����򮠠�$������YV���W+�R����_��TUk>{�K�3z�U0�`�ڧ��6�f~�a�˾A$�W)��\T=������U���'�jc'L���]7V�A���}� ��%ր����`!V�h[���_�dq���Fɜ���z�r'��B�R�4�>�
��W3�1p#?�\W���rX��8h���P&�?��^K�����~�K?�7h|����D�nd�8��?e�cOR0#��2�����k�B�+�G{�uc���CJJI��	������������Z��>x�e�Qڕ��g�SOa��X6J���;����K,�9<���ҍ�߈b�x�������'(��ƷŁD���������T�mD��>){[�L����������w��{��&�F�/��R�;ż�iu�k�&����߉%;�w�siǮ�^�}Y��޹�}K+\��T2J ��IsU0ݴ9}v���e�fO����T��3+��Q=��X�0�2��5.� 6��Y�ҸM��q+� 7�*o�T���<Q�+�;e����`��?u��?L0�v�ػI��b�zy�dqu��C�%�.��>�/	=~'�T�6x[ǐKB�KU��Sv����[�q)�nzo����K|��m�8����R�`�̔��:` 1��I� V>�P�ȥ���:�| �d���Q1Z�2�u�2T�,99�,�-��l`��t*�"���t��~r���V��D���?Y2�:�^3��q��aQ]�I�Uy�?�F�{q���wl-�_s>:��V�_u����ڗ�0-�gϤ�u\&�(q87���R�H�rv~dd�?D�WJ�D�I~��΂�O� h�>�T�$uU�6�x�	/���� G-U��$�R~��z����<e����򹌆�
Z�'�n7�b5޿x�ٰS�@@��&m(AH�r [�{�� �3�9E!����B�E�_�1�wޑ���Β+r�8��`}tR7��͐v���`�o��Ԁ��t���G����tRi�8�#�(����t��ژ�J��')��.���:�
qzwy!q9z?o��C���O��'������D9�������>�����r�����T��Df�G:���s鹒ᱺ̱�Ci.���=H����xT^4�����,s..���-�k[%7�Vs��џ��L��ߕ�� �������t����6��HN��T��$�V�v�]o�ǡEX�#�R�]/0��GKMET�CV8�^�)|���|X��^�����xA��~G֣D�&� �.p��t	_�f؂��WVA�^���Є+�K�ܖU�i;^ի�1QSS_��P���#^��
e�_�jh�W0������l�z�`�h,+N'QV���V���';�n0����l
��~�f��V�#+r��3i�g��m�_�?L(��T�`�]t�j|/K�����z����r�Y���eF��f�l�gJ(����6�;;'gs��[�W;	4.�[7D�6�|���X����8zI�AȐ^���qo�N#���ys�ٞ�MT�퓿�x�C�xi@��ôz޽����ф��Q�X�Yէ�<J����F�?�����*�����j��W����Qɏj@O�p�
�	�\}1f��Q8�Q�r��ǩ���דy�)o�C�-�3�u��A�U��ؑRWO�e����č_�>��M�Pz�-w���ޕR��N�Z����Q�^�x�Xkֵ�|�]ҭ���,;/(y�+��������,������(�N��6�6�_��ɏY�eNI{���ֹ�+�(��y"l*l�"W5���$�fy�s��[��m�}��xA�����x¼��唶l��k�׹?;���+T����N>5��%���)O�l��g;F��5�x�u����[݋F�ͺ�	�T
�D˲m��uu_�wn&�QG�˅Gu�\�q���b���M���j'1��܁�YK��ҩ��'a�^��^G3.����������r��������A���2���eWq3F�/j@�V�����!�Q�^�����9	XA���QO?�-����X��bZ���U-��r�?.��{�=]f�)���sn^��k۫EGr&���M��<6l�4��kW)3+���ڇ��4�r�6��b��}� �;lY�yݻ���<�^T��^TkVҝG9:!bVL�?��V�-��K��v�`�ԍ��ŉ7)��}6i�J�@>�]5��c4�ː5���tw%fx�JD ��0BXb�N����V�I5tka���'ğ��\C�RG��ϡ�G��0�����/�[b��K����	'��\�R�����������D�,q��l�7o<C�3:+�X����2=�`�-��Gu��|��Pvx��t��(���x�]������⧟¾�4�J��|2��Y�o���T�#��/cK�?qy�s{�mA~�i���q�i{�;I�t�ƀGAn���>nE�����仩�o?��xM14�R�*ȽI�K��|V?U:.��O��8��3?k�}9�X�r�ܡ��K�t�?[�h�U>�~�bp�i�Q܇z�rq���n_��:B�G�M� ��=�B�&�b��f��.����QCp�G�Rr����@UC`�䶖�k)�KwJ3&sa�X3�]_z�y/$��7m�R��2�jd�)h���Ae��(~q̐=�w���|����پ� 0���a!��I���O�,t�j��SQsHTO�����E����|#g��1|=��������?UԱF�6,�x��|V��5�oWď�+�N{C�O ��"""��3��G�vI,\zO<�\��~N����+6����_����N�R*Gm&ښTJxtp�0�����������ALej��4��\��N�Vo���鄚�r\��fC�--�~�ao!m�u�m���JK[��� ���q���iJ�,���?�3<`rtr@⣗�C~[ZZJ ��W�V����&�u卦8���!���Z��@~L�[�]�;b�s4���n��ė0b��������NU�_r�8�+1����Q��\�5��X�kUp2���"�m�{b>�V"������p4k�?t��B�P��+դ�Dt�4n��`���(�Л��Q*Ȧ��ײ�A	\��p�@�������W�<���w�4���ͽ֌Pb�G��������S@$����k�垺K�u��[}Ɲ�i�&�u�3?������'����(��
�z~BOAZK�[)�"J��[xL��I���s�,i ������������T�����<U�ҋ��Ї��V����dϐ*r��&4;;�junD����Ld8\�jPB���v�A�+���u"|hA��gE������7Aao1�>Z��!�+>����L�f/)K�=v�!�AJ��O���,�W�p�T����`SV�b�R
�_>l�f�{��'?5M� i�����_�Ik��+�B9:����3�1���<�$8\�������=X�ͯ�����P�-�m�W-�D�6��@�g�<���𖯺c����?G�,��?%���V�"{Ž6̺#rQ��yq����(S�Χpé_bO4g����*OlC"8c��Q���!�j��;��1E��*��\h���[5B����L
�{���e��а�I���˾�*j���(:O�7�,��I*�{*�R �d����͏r��R�nk�e����4����	��QX�=�E{U��7��j��.��'����@/ؙ�K�Լk�"E��Z��
�;�G"w0�}1�0h�:V:!�a���c�_�&����cep�8��՛���2kh�[]___�T�a�Q�N��bl� ���h���i�q�о�m�:1��d��k�����[/2ֿ�`\���+�A��A(�M~�
D��j������
.��O��e�����Ԋ.8w��睇�!Q`�g/���ppe�G6����F[��6������m�6�Q��Pg�:��o==T$s��ML��.g�½!�7�:�	�M+x訾'oUxk�N���I�".�/O'm	ǣ��m��=�
_�]Ѫ�{o1�+H�~�V�Yո�[��z�:8��
���:�-�}[���+M�s�ᣛ��i*G�˓�;��Z�%w�����Y�-3'��~8 ���J��0\��ڞ�E�&� �KNu�8b"�����ٻj����eK�"��yߑ��;4�{�w�?�v�����684�F�q�9�e_v(<&��>�B����IY̛!p5<,��,˳i�=�#��o|{4 ��ZAu�jbw��N��$�����^�����G�T��h{�1	���I�UXt���G3:�Zj�[[���ђQ�cM^_�QTZ���TT�����j룇&-ˎ����{��U�ؕ-;����m�d�7��W��F�.��UA��.��͑�� ��D\ϾƠ�[:5=���  �Α��`e��w� ��C�o?zI�P��M�r�[��D��˦�۳�$��8w���Y���n@_h�rXIԓ�έ;ƃ��w26c�Ėdܤ������Q�+��Ӫ���_�D���-o��>� ���t������&.��``?��-�h�Zb��s-CԀ$�X:\��P'�\����#�|����D��)��zz�SU���j� ��`��t��i_���LF����8�G����߯q�s�;r�^yNP�ӸR� ���q��z�����mm<c��,_�Q����c�F{����y_>(�s�<����l̎'j����TҸ���&#>�a�I���C��^��~����r:S����[ uL��~A`F��		�z��7���U�Ŧg��7K��PP�����f��H�q�j��I@m
{�1���ۍ1���X���&�q�϶�$1��j���L�
������J���Ι��by0B[n��&��>�,�E"�>�4ݙ�6GCwg�tXϲ
�)=xÙ �X�e�Vt�����1�Kךm@��:�xVv.ޛ�#����������D�v�W[6� ?pj�%�v6.��žVdzS^s{�8�𫨷)�ŀ��);����Vt{ښe��e�W��T_1�,�D�Iɳ]ץ<�}�z�����1;��¦�T^u�C���w����J(|_n;���B����F�n�j����đC<�>)���G�u�W&#�2qlT��:
�ꁷ��\ݦu �kB��ҋ���q���mQf'��ٔ�'�5`�/�3��Հ�1����kx>'�����5���;0v¹]|��<�/&U��}�۶��:���]�������0�A�������y]�_���,G�=����D���6�����d�A�55u��B���Ə�+����m>|�pitq��cؚ]���1���GH�y���ε5���<�=E-�;�|���\��yb&��N�����tS��:�ӡa^\ǫy���[�9@�#}7�¶')��:���1��&�\�}z(*&����Q��\ɾ���cd�s&I���\ӯ� ��w�����&1��^y��;Ys��v=ֈ�ҹJH���?������F}��]Ϟ=�c�%a�I��FvvN%x`����ҭ��1p>wSVO��{Uu=�u!�Սj���%������iP���_��bjZls�B��(.G0�.�zU-Yx����{"r����]�Vlv0VN��y4����d^D5V�8�&���hz��tѵ"�c�_��c��
<���\8�4�>��3b������%OU���kmi����.�?�r�d�&���@6V]gy���v��g��F�~��@����l���V"�)4��gt�qoHws�D�i�L{�TM���#:�ڼo�ρ��z	lJ�[_熽h��7SݩҗSE�Ӥ�wf����[��x~���v��9�P^�`}S�jZ�hD�i���JF�E�C^����٤�����h^����*K�q[e^+v��߷E�!V֋���߸?NW��f�G�W�7q��gg\�dK���9��W���v�u�^׆�~�2�^c���OW�M3�lM�m�(�
�P�V64��E|r8􊮘��!��E�΍_K)L���b	�Xn���f����?#U5�Q11�"iR&%r%��>�,�m�nF�ش=sI��y{P�������CR���{ͨߒ�1/���P������8�j�G�k.�� �2;�U8���;nw��z������'��1�aP�P���#����)�kn���$>��(�rk%�r�鋆(�>}��5וL�3wV���;{�/c`�֥����� A-�{�ޛ~���ٕ��	��8���������ɔ� �[�qq�������^�;�m@�K⧭xK	j7`��q�\w�r�q��)Ks�-�Z���a1ٝӜޤf;7i������\�M��ĩ̴�L����q9o���6�m�<i}��_pSS���b���Y��~�'e7=w���^)y�ߜT;��h���
R&�=�/�d���D���߁�%�g#����F�T�������V��k�m2D�%�fQ�_%���m:s]ù��K��)����zzzU[�?GG��#Nwu"�,G�{6�O�{�� T�j9|������y>�ϔO�&�!�o榇�7��E�(5 ��Yvw��@���I��;_58vb�]F^�l\F��2��Y���@��d[�{�'3��i�un���M׎�r(�֬�w2N�^U�=�n0ڦ&3-������1KGҟݹ�.��N��1���/�2c����=b�o�S.�|pa _U�����J���՛͵}��]S�g�|7ȏ��7���1�T�������m��ӯ_n^�����x����5����ޣ<~��7��칺ۿ�>��m��u�����ډ��7�1�d掫g<2`�KI.�U�y�z�T֫����`�?������;���ƪPBS���	.X���5��$��5G�fƭ,����@���0�i��h��T��ȕ�b�j���p{�2ngLy�1G q��	�^�P}�|f���J�:�j��qX������*R�Y�K	��r�[R�<>���"M��a�O\��Q/'/�R�����Kq'e�4>s ]D���-���3119�X�W��37��l�rX\⋀����ܞ�KߩJ�蕭4s&UHz�]AR"�/l�`ط������çR=.c�ymmm����i]c��M��珛�9��wq�=�p�%%�B��8�<��2O�� h��]�`.�<P^��,�ţ�W���H�ұϴ�l=�]�a{��S���sx!���IZ�7(����������#/CKf���K��-�k�~(��8{A�H|]Q>�:�RTCV���Xq�,O]511������̲�������.�Wn�	Q��v��G���h$�\F�h�=ijj�z`�|W]]=U�fz�>6���W�!\ⓣ�OAN���bf||jT79���-�C�d ������]7��Iu+����:�vX�"��>�B�����1�)�h�����|�ΝS@l��Ċ�G���i@�������mQ��Tju#��4x���P4�4�:�K=��0mV���u����M�z��?Hdk���l-�,��eKe1K��ҁ߫l�Z���� UD<�&lߍ`L��,u -Ҍq�Q����	�TaS��ȫJ��=�?�_�,��f�����a�dWkv�ڎ�A���ч t'n�9ȜR^i>z��(�Y!uԀ�n�$�`mr�J��gl����I�X��f �}��H¤|�p�����^\��g�K���!��k�/�\��L���Xb�_2 ���]ȨϽ�̴9���@}�w��M.133�;!6XX��C��Dk5L�!�ԯ3H.G.��l[2�/�2p5��D��U�VەURV.�,B���1����'O�e_����L���Z7ZG8��p[饐�����Z���t�lF���O/W��0S��v|!.S�1���E�!L�d��Ɏ�<Wh��kk�����w`;'���K�Ye`�?��D&f�e�	.��Q��@w�/1���,OE�W�JW�!�-g'O�<U?����;]f�K"��CH�uׅ��h}�=i��l����V��.�x�[8��۽��e�.�D������%��� ����}Z�-���2�4�B����|��j�`�Օߕ��g���>|h83�Q�2����ٰ��v���꧹��jr=��J0��R�l�������/--=���6y�|�JfVV����r����W�x��Ek!�����?EN>�ʞY�fe������}�V��d��7]�tؤ�G�N�ɠ�N�?���2�nI��ޣ>S�dd|=�pu�z�����5���}���O�uu�jjj:���,��vU��E�$����'������#�$�������x{jû|��o���f+�p��:���,5�����s�MA,"��w��_�}w�����d	�S��}�w.�=���l�H�Z&"�����d�~���}������%�:y�B���~0�y��(tL\�qZ^Y�x8"�E�!�~��,�(Y�o�cn:	u՗��Td�nmI,���57�����9{x���Q������EB����˟�����(8[�[��A�豱��|�)�� V�����AEN���,?���O ����=�8�&�4�ɞ~�:8���qΊ��cà��i��[���,xg.��x)n�����%�}ڵֵ<u�r�;�WJ��`��l�Z*��"�$�����3S�΂�#�F����̬ �־~\�JKf�k�w�����p��p=?Ԅ�#���O�Q�M)��h���#��"�=׈~�N�|������V��d�lg����*���ٿ�f�_�;�Lm���v���A<	�����uz(�M�W��$�T��o�o����#�55q{p�Ş�k���ZG�@%����!��,w� �
��� ��a]����H����)���T^{,2���������m6.����l���#�SZ�M��0?;������۽8�=i	��"ps;���g;:R�����!԰( �W緁�1��oTH����Q?�|V[�x�ؾ�C�;���CEM�GA���3G�>���CD���ڹ��ǚ��1�"�����U$���we0�+!�ّ��HnTG����O�\�u����]��;�����Ilf/���@T���_rAt*�d�X7u�8�P�1{�r"���҃|�+k��l��\���EMd1��C���������ײ�rt<:�TwZ��B΄�Uq�IڠL窈��(�t)�:/Z�j�pJ9��j��ׂ�¬������K��b5��VxE'#r����84�5���]�L��Q���4Il�p9󅊓Y��T9��w�����t�)�#m��;�;<&�L%|xH�����Cv&)I�mv�gjXa7]��1=��#�l�±o7� �sX��&M���C�ޑx��c��WY��5�ޏR�7m%id��
�!�_kVA�4׉��,��]�u�R�@{�I���x����8,lI~9z��^]qp�$�ͣ���78o�����d����g��Pj�
�K�D�}pg� ��X�"�lr�"_Ѣm�韴T#d��KA/fI�.�|6&Ue�r��%.�T�Ti s�C!���w��t�>�x� ^f��
XK����.'��ܢN��Ng����%��r��n��G����O�U�u��Ύ���e��|�JUg���gz�:����l@����ظx4�:�u��%yB�!.�R��J��T���
�%p�w���e  �i��(Պ�CS$������U�Wu(jn�oܨB�5����Г#�	+�k�������P��wo�(��)��d�jW�x�?�[�6���=cZ
!���F8}��H�=���TO�'$2�z���*����?�VA��@h�C���c@�{oRܝL�۲[�<L��[�譊��E �VL��Up͡� ���d�RS��*#�>@�o"8�t_��1���_�wxr{�@���GY-E�N`j9����N�|��_����Bk���A$t|�j���v���W"�2N��sﭏ��{l��|Drܛ7oznL6�~��:p݌�����A���^J=�;w����+*&�z��f܇���i�����QI�r=(�3�#}Mxؕ���$eh��(����fQ�,��%�ث.�Ш�,��=~�AW���B!�{Y��)k6_<Α��[�ML<�oʿ��ɓ<����	c��>k��m"�KLL�M9H�1��r��P��/X��?2��mq��_�/T0���������WS��i�Ke)_T�X�� o{�.�"�>�Uz�T�U��x��i������#|�N�<���w��{w���8���e�b��pA�.3[���h�����j�k�F14F	 �4;+�<�ya�cV|�%�$N�!Hq�լ>r1��#G�J@ȵﮡ�w��l"B%��^��W*��P�z1Dqt�>F�[����/pT�_���n]B^ N��1!�T	�1R5bbD~-�ލ��j���Ji�Ԟ���C��KX7��"��<�[$���XZ����z�����ݽ�x���vu}*����h,�u����+b���aϸH�i��A;�|R@AO����z��|��O.�ǀ���
��N���N*8�/�����ܔ��}�/�؏�y�n�E.[v�M:,�&���`k�m�k��K���T8�'W����62q�Բ���tB��]���^��>��I�(HT{i�aib����Kc'�Ͻ����j��c��i�<��A���ҷ���ڌ�_�``�_+̻�d.^�1n;� �m��q����TC�,�k&,"��u�������ǒ�`j�5L���[�$ p�^�,Q��
�b�{�F7:ÄVG�_�ɴe0����x���d.��]W�f�#�2��;���,�$.'����@g;�q-��cء��2yڕ���#KgR7�����&�)�%u/���(S�{Lv����l.��y"��T�o���8�x���MpPA29Q��M��>K�����'��u���O	�K@��
}�;~V.�*@>���G����u�'bY��zC��.϶"�(��+M���B{"w^��V�A���KR��)\�ŉ�w�s>��+�.�n|�nBE��'5ϸ�D���8d��a(��IC�|5@��:G���C��.�O䟬�	=1b�Z�0��' �B��s�wԧ�{�����"#����%���qe�q d_4���g��m ���׏��޲R	�)C1�1_��f���r:;;z����U��%>?��zL�bD��h���bMLLd[���3��;�P{���8��<}�����R� \��`���c2�:��?�4�"ʽ�Bt������u_�3���w��ܛ����xo�*��m�WI`�����ﾸ����W?��X�Y(Y���e@/��yo��S�����vޤ�� ���8�q2��-��=����t篡;ھ.G2��u�o�'�>qr.����k�	ۚ�e�ݵK�s�6yް����%�� }E��ؚ�se)Q��~Y��<ʟ/��/o����5^C?�����E��~sc\�=�dt���5��}-p[������(���]�d��A��<,���W}��xh��q�4��]�aF�y�<�|�"�́!�c?����1	�ac���MGfq$�7
D���-�,�W���jk_!Z�a��p��}�˓=;d��W3N�����9����v{Y!3ߢȸp(�:<��\�|�ߺ�"i�&?�zo����z�i3�WXޤ��U�:��-gj27	�s��
5N���ͺuX���ҲM��r-��
BRv��Vʉl,�6��&�����>�У+��̼?ނ&�`#>�؟���||���x�ΐK�U�6��ߨ���T��U�y�m����郘E�&b��3�����qi�e�������_�s�c�>5���>�x�G�i���|AҒ*ш�}�M���ܣ��YA�*�9z�h$��
6�QO��P�s�=xF;�)�ؽ��D�5�{��������P�ˠk��P�;RO��b��=��[���Y|@*+��?�AG��ׇ� '26b��S�znF������A��:MC�ȗ��2'���9���J�繋��1�.aKo�^;Gڋ���șF71ӑ&���'$���W���|�����h�7�coM(�p�[��H��W	=���i�g}�C��D�O�������v�'e���s�jTLw�ܴ�<+�G�E�1,�A^�=O�߂�^"�MV�?�7�&��.Ad \���/�$��Q�eD�s��&s�#8;�0!�V嗫b�e��p��Sz�ެ���)��L�ʋ���wz�=�T������U1�6w{y�]Z���d�n��D��g�r0{����?k�q��ۄW��Y~ N����О�Xu�n��i��	oIy��r�.����/�^<=~��+A�J�_�	�����{�G0�'����۴j\��3��6O�$����& ��Z�7p�,����1��2���9�Jq�7*[���� uѷ	s�R�|D����M�1O~t� ��<� M/�w�+�&=�!�ܽ�|5�7��J�a~�������\���<�p����m�,������fy�ٗ��$k�h���D�[����4��������$C<�UO����m@�u���u}t�<�e�����"�Z	7~xm/0S��c�@��&܍�B�<���%�.�p�?����"�A7�9��m�:ٹl����C���te�4hkA�����2�jw�����)�f�����ku����&�l0� d{�����se�wy(�����m6�v.��.��l3��v<FkN4==�>���� ��9셍���b��h�n��/���q--�|�r�D�â��z�D�q5�0c�d��/�<�K�*���ᴩ4�8�"���@XcA�<p�3C���0��3iqx�IsE�g�A�#�ר���(�i���S��������g���I�1��m��A�_�`�klJ�㦌K�l��70�Y�h1�X2���^ƬX]��=�5d$3j�0c���hӿ��ၽ=�"�C��C�h�h�	Ԭ:���嘣KKKe���g�O#l�.�����SR0 0��g�Я�l��LRg��(yˮcH����,F��i���Z�q��;d�b����<����n���s�ܡ&PP�8�F=��k��o��p2{��]�E]��	�����G7 (1��{i6���_:X�'��䙥�u/�#x`��z�߇o��W������~�;�Rjz|�ֲJR���((-YS�e� b�]�*��/�Ik�n��j8����^���14:Q룜�� ���Ǫ�N���������b,]�1,��#����yӊ5�}_���U���3�K��?S�j	���Ls:"�y�0 nk�E��܂��X�T� o���P�7��p�a�T�SN��N��=�>�Vf4|4a�����L���&��J�86��%�8�)�I���-���y���<��֤�i�0�Y��@��^����u���2��8�<��x��)�rD���e��.�`t���\�$ڏ��T[8�^������7�V3첽������ruNZ:����CM���[�[���cEi&h�"�wê����R�@��uh1�a���7��\p��묢�;&<����G[�W���9ý�u�����d|!]��i꺹r��YGiN��^.�������[,���|<�ɵ���e)��V>��u�v��_��W�GQ�3E���r�
���d9����m�N��n�z����z48v!�}Te�pB���D��=�z2{'P�*R0����B�.JݺAUa�3?�V��
������DP�[��^g��X:�ΰĢ�Mzu�/��ͳ�G߅Xb�V-�UC8Ƥ�#eoOSqkR�1˻��X�?������5���<4�l���v�4��b�'� tvnn��RȜ*�7;܇Q]��~� �b����䛰5;�
�����x~��l$t�T���$��5��坖uI���@'Q:����l�ʴv�_�ت�.0�f�j�@^�o�m�.$<}��%��y�Ȩi�T&!���-�J@սT�D���I
�FL�T7+��'�-ɽoU��F�樨G$ O))�=��~/$Z1hM`������D��P�����2����4���;p�[��{�g����A>1�=i��ۉ7�iFL9�C!���̞Yj�P�5e��L�F�������-���Pn�Nx�GL0���}��5L+mn����x|íb��;K�D2�Ġ�p������F_�Ah��'w_�����Z�T;�������,�8X�,�>p�iY���7n�i�/7??@�t�a*!�P!5�p�׼Bs��?��s�jNf�ϕ�� ��Ƈ�9��X�� L0�J�6�F�����rmu׉g~��"�7R(���nhDۑ/g���dH�@�)#H�;���k݉��_U(����n��'M]��a����]^��'_��R�M��#������]t}��aC�hzz c?
�_�wXH^�.�ዂ_�9��D.l�J@>�/�}ت�V�4L�U�=j3$��&T��,t�ѹ�o���[9֝.��/w�U;�v��s�b=8[�♜7��Q?V	��W�U�Y�ZP�x|��������������?��q�����>��Nc9q����sݜj����IU󳊆�D��	�]eQ6�,x��6fLc�j4�/i |>ln���D�aؒ�l�����J��1a�Tˀ�����Y�*Θ�ʾ��m�^Jhh���H�詈�d�j��O�����R��K��g"h���s;�i0}��u���>z�W�*�H�Ɲ'����h�s�o?����^��@*�%�E�{_��mddem}�&�o���4���YW_*�<iP�v�+���o�"Eg�)E���M����KY�=��?��R&�4"}d{�����7��V��c���(��K�������l2���d'g\* ���)mU�Z ~�����VA����;�Ʌ;3#��
�s��&�����\t� �q��Ș-PX�|���ѝ"��ՙ5�ض��ԟ��%N�뜞|� �u�x���D�d�����Go������	�������{�����5*bz8�eb���R"�0ziQu�����0�Q��b��H�͓�������.��k]u��ǝu�KW���]f~����Έa��tI�fq�'��/+����&����q�44�׳z' ��mUf����0W���!�z[
�H̙��.w��d\���#�>���JJO��xlO���Z\��cߞL𤐽{����W����f���(^ߚ�<��vH-/+���$��n���[�la{�o��{���%r�OY�?�v|�F�?I{�B�;~ ���[ѭ�q��&�4�o��YjF���g��S�r���Z�$��P�2�Շ8Xji��1IvĿ��67Q�t��ͻ6���͓D����V��ǭ;��E4�S.ww�i��?,�Xv�V�*0em���uu�'��}��*� E��!Y�N$X�#+:�=�F0D�K@r�I�Qr�#���pw|K@�Ge�����x�����(!��E�M�3D*#YWF��q�k${��ɾ�.�ȺHH��^��6���5��V����xxؗ�=�s��u��uYm��A�|jt����D~��ƛ����ƃ�\~�'�|JP5��6s�����7��Z�/ �d��]8���9!H����i�'����)ke���	N��y�_r�&�6�֭�mD��zд���=P���\�ᾱ���ǈ�P�ڥ'a��ͭ�`D�_�4#7g<�i��?`-��}a5��>�YO@7����<\���3lMm��`��S���*��IZ�6��8����W��ԉ�l?�	�^g�Ҫ�V�����H�ݙ��sÅZ𑉷1�S�
6���}<����O���R9����FJX;��L����bV��ٚ:�/xM�������M�|t"{���gb&S���te�Ѯ�P��������	B��,a%���<��)Hp@���~<���u�����NR$g���n :��4���bT햹�2�+5�'��~/�d��~��E��
ka�Z">�[����3z)��:ŪkgG�Q�-<�J^]ݽ0*��,��w�����q?b������}ݣ�[�nǾ݆i
j�J��+�%7ا�����Qv0�~~��+Z$j�p,����H�}�zs ���p��f�K����޽E���cF�{"���?�>�\�?C��5�X'�%Fl*���7>|�A�*��ھ�G���������O����Y�:N�i��;o�4�F;@IJ��򒪊	��s�
��	��z����y������״�e��h���f��FFc�N_���fV�~l�me'<���Q�qs�JE�༎x�[ )�1,����ZgbW;U^�1V�Q��H��8�S%�i*|�'�����eC�G�P�p�5�?��Tz��-:6L�UT�;	S�;�۱��)���=�D@�ږ�`���n�-����ȁ-8�:�܋u���~U{s�k�����NA����V'\�U�w�uL%�yLF+ϋg!"q���7�Ŀ�0E��U��uߴ�}��염���vOZ\@o���~�ư6����r9�HzT���k��9����D�I�N�34��-���8��N��NDT���HT9@��&�+ۋ�̧|���Z�H`ܓ�#���-���x
-�b��D�I`�6��{�B	�K����I�3�����^`)-8t����6(�E%�29y�OD������U5�~*RI�RG�	�w�6�$=�&2x�pKp�ޙ�24r8eLz��5�U3Myp�x���x�g�������F�B`�Sr��Iu=�fE�ӗ�I�'�����>���� ��9IK�g��y��6̜b<ot14xϘ��C�[ �Jbr[j`���S9�ן8\�aY�Nֿ�;j���[ ��=�\,�>kx'QtZ������|�;�u�
�R;~�Xo�[����K�"p��b8KMH<���)�K�����|����%���+�Gx.�&�����������zߑ�D�n��`0;���{э�?���F�TLY�_׈�v���>`y�W�������N��:3��/D�7U�_�n[b��zj�RA�g�F�����~���]�)�ϵ��*	l�da~an��7�hTy��^�g6����2xn˸
'im�����a'i���3g�e���`��͖U����$�((ɠ�r��S���U	.ٯA�b�6g����/8�9|���ǫ��n�%�7��9s;�u����V5cj�~��$��R�3B�V8���{�éhu������c�掤O�=��~��o]&�p�'�:H�{�ǡCM�IF?�0u�>]�����47�mG[ݎ��^k�>�UJ�������+ˋ�mǢ��z��q����oC�����v���jfEܽ�+�=���|�у��^��_#z��ܚl�Q��Ͽ���x
9^��� �^����V��gNI	w��ಌ�3�NDssW������2(k��� �i}���_�sC0r���y��� �d��~�5*���1i~�+u0������ s�ݴ=1��u]�z_�OD�s�Q0�y��n����ln��e܊�t���zI�#�~�$�k�g>�� t��ڂ�P9�J~�́Ć�h�2��lFcS������&��c[��.�G�Y��z⹀�Ŏ;�k ���o.�� �l�-�(��d�Q�y�ȕ���7Y�1;�:+&���k�"�V���z{�T�hJ��,{Ȓ�F��1i�,I��Z�~����0tmn��H�T�QϠ�2������e^�m}��V�B3�#�r�1$i�ۡ�=C,!Α���ځ��p���7���ƛT�S0�XS�����*} "���f1j����=@zA��p�P�������:�ܼ6����}VW�ɲR�S�u8r�7/f
���M�	Y�Z�B�ùT۸�C�~�%�Uܙ
���ݾV�v*�l\��G���?U_n����pV�]�LW��y�p�6�y�3��TGֳغ�������}V'�b�=������ ے^��vV���q���F�9\=]��Ǜ���:��*�m!턶u�m`\x�^�s�J��k
}Ѵ�Vɹ����>Ҹe>fW�t/��6`��^U77+�z�DMMmKH� Q���)�n��2m/_;�?��Ư�hٴ�zr���f���嚪��6fe�c	������c9}�O���d������	��P�1�B�U��Л9�Vg�����*  ��K�k�����BTTT_p�'�+�R���+~���+�>�Z���~�*..�/۱��m��-,�L�"��z
�D�5ɪ�h5 _q�+//?�����N�ş��̍gc,�认��CwQrq�q��Q���)�t[��)nf����f2���3^��m��UNp*|�^?��qb�CÛ5g��.���i�c��"~ Bt\��B�I�Ґ��V�_��u�֚j���Ό6�)�W��Ln%j�/%DEC�v��n�͐F���$�.����}sf\b����
3�9�[R���5A����$���GMVI�N���-+�B
�S8y'NNI��z�
<�p�����-���?�N��S9�v��uf�D�;lλ�o5�7�R=~5��
?gH-�8BM�qs�Ip�-����v��Ru�Q���cdB�A os��5]��ocI^7�Zgٞ��V�=��S��:����˛�Ξ�}��+����2$�#�gK�m�~��U��2�J��GU�0��:�����J]����M�2�<��؄�G)���Š��3ζ���BWשX���l�m�=�2=$�K��������@?�V?�m��~Rv�{'B'm�9؜i�!sn�@0U8p�dacc#�B�É*�����l̧	�}����������ߗX6�
�^�����1�R����#�W�9���`��Q��>�=#*��X�c>�x�����b+��E�+�<�:�<0���@;�ug�*��싞�����l�:\[��h�8�d��v�K7t�<\�A>��i6d��q��$]Ӻ�s������J*ԋ���ܹ��d�=]���.�jv,��%]sY����C������q��B�l	���sQ�K�9ʹ%.<u��������Qr��4)B�v��=���n+{��&��2��7m�L�m�3b�ʶń"�E������Sљ��AZZ����z�ӊ����DYTLlع��׌��羅������!c�Y��������jDsHp�:a|����8�������RX��y��́�'Y��Y#'�"?��͔��4�*��x��6݆�I���RYYy���8�tB�����M��v5rI�4��yi��7�_f,y_�/<}Qy�
շ��j�`�׈�/�{��s��9R&{�g]��t)�W&�ʎ
U<@tF�Z�o�4e�!�����nK ��e*_���8�(#���*N<_5S�����g��|����X����G���r��*!^n~O��/�iw���T�'���2�e�pu�fU8��7c�Z��S���=�O��!	��E�S~e �j�͎�OZ�w*���vǣY�=�Y��	Wם��f����IZ�1K�A۪���;�n���Dz���e��ñ[��c����Ӻ� ֺ���S���ӷs�(�3���*߾�da�]�m|�,U����CzfNM�hN���=$�8�{��rȵ��u?�s�z�����B�rӕ��H{�y�VPљ�洵�32�!FGS[  ��H9Q����	ݙ�i����g9��������@v�l�����J�v{�\f��k�.����,,���ݲK��6��8OЁJR�*����2���b;+ߥ���u���=G�Éҕ��m�����RY	��fj��G�~n�z�:��DY	�@g�T�b������[	㑟�nm�\�8|��ƙ��On�Vf��x�d�c�v�oL�b�J�S� )=n�R<e����.η����1�k�34:��m�;���S�vf������#+���e&)�E���ǲΩ[���0�z4���	|��^�_/=i^1�Xvd��c{=����|���l����腶S���ں�Ku�����N��>uW N]%c���7�6��/IS,�.'-��Â'�� �k��1pI�6UG����vO	
���J}�5��_w꽿�� �6/��;e�5�8��ƿ�K2��"��XU��e]8�:Q�xM��'����jZ�jh��j�&D��K���S���G�SAx+� �kڔ�����c8��õ� ��yk\+�[�(�3����N/g�7����%ܖ%c�Wm'�w)�%�g�Bv0����P)W2�nc��Ґ�]wrDFޓD��҃R�h,�C��g���:��O������i��B�,g�be�ј�ũ��6.3T���׉ �M�%�_����<��+��qJ��zR���y�'?�G���E9~��բ��U�cK����������Z)�=I�p*�EX��P�cojaV��M�*�#cD��&"2퍹?M��Vt�aʭ���4�o=����Խ<��C��&s�Ȣ�5�����j�p*����/�b����g�#Rq։���$o�����6���Z $O�S��:�hy_%%�� �~�B	���XP����Tu�v��V<����LIu�]�e�{k�����;��Z�	������1��R��|x���3_I�1���[j^����6����8�*���-���_�2t��[��z���o�@8g�ž��C�8�RܪSe��RK�r��M�S\���qK4��������MJ=�T�+v|�Mj=�b��~#����� ���Wn��hH�H�ib�B0�G>�ͩ�,1v�����b/���߹������J��/$��S��Ho#�7���ܵ��_(�e1P�c_z���+CZ�m�(SO!�lz�rЮ���d ����<����_�`J���N�0/O/}�T�Dv�h4�;z�>�a�"�\/H����jk�}I�w��Χ) ��v��{�6��4�Ѿ��Ѷ-&U�٭-q��tBv&\��b��Bi=�P��5x�[�F�	Ug�<o|z�b&�9��C�Y��G�q�n�|� 7���6]�El�סw�c�r�ǯ -�L��9q�;Y��۝�;<�}���6���Tn��f�M�)E��1�7
��tk6���:�Qɷ ���^�w�#�*����Wk��qK� C��9L�I�=齾��W��s��(~��ĩ���>�zrL�[V �e�㥒t�	N�gcN k���R�#��Eס\L�R���A�����fkv��\%��3>�8�KwbA�Q{���}���_n~~1�cRP�A$�.��Ս�RbЉ�:&�e�\�\�o�x�X��>���K�JH�!�}��Dj��+��������+�6ޝ�{g�s5&N��s�0cf(���hI��0�v�P��]!����I��U��N�vtU+*��P�R}�W9~7 ���XΤ9Tp=!���*Z�/���:����E��U��k3q������6^=�'Rʥ����iQ��<��f�V[�WZ�N���y<��p�:�u5��s��,wy!�f�Yb(H�!o��"͐]��r.q(W�M���5u��D�;�����ۻ���r.�n:Av/�ĺ�,Y�*-����I?9����m�J/�Gu��+VRm���=Hs�R����S���t�u��U�?��^�af��J�c{��:��8	TC{��C��u���#q�Y�'���g����E�~��_�SsM���C�iB�v��2�$�c	�����V�/<���`f��[��E�l�^�����d��H1�Q��aN��-F�X�hoE:�\�Zw��wc���6���'��ϧsm碃<��'�o�GM>J�>�#c�;�����c��DRH��/~����T.���%���M�v@�R�.O�Ӓ�`��cn����'M�S��ͧxm?f�F���/
�*�=�-ڂ��z�@ϩ$x�O������k��0_��z�����x8Ŝ���z;��R��� ��/;�@s��F^d�2;��:=���ykn�@.F�r �Sٚ����,mx�C7o���әtz�t9dc�%�3&�����)u��|����.�@����ka�#���^��s+�B�mc}�54�.��/7�r*�9܎�Y@��<	J����[7��pt���Euk�=6�:�%���������R��8OC#FP|���vqc�y�?!O�ڪ�@mԭm;#��*�E`��oOW����Rd\�./;�y>���zE��)�{<	�X�"-��n�"M��5�#�@��R5ᠩ�	�[X�&�3�Q�����H��"�Ӓ�I�j���M��~���%d� ����Y�(������ ��>��;Y@��lY���C���g�s{���Ar��H��c���Q�l4r
� �D$��}�]K�yʺI���m|��o��g�����S�������߁R�.��{�rP�]������~�y�������4�ב ��ڊ�l�4َQ�i��P�q�Mx��T��QJ�淇�zƱ��yV�
*W��'�Ķ�p�xy�mf�So��x[�l��������ކP�6�!�-�þ�P�AIP�� ���~�����!#M�џ�T�d�T�T��|�뎫��8%ů<��/��%�F̪�[��f����禔M�X�>�z5j����׍�v?[�����p��}Mp�U��F	��,S����m�Ej;�-G��n����������pD#����o�� |t��]X�D2޴]ІK�����O�4G΅�S���~�H�����+S�føĠ���:�緅d:�$�|�8���H���p"����3ox���%�<�s���Rc�ܞ�Q֯�boq�*�Og@��UM�F��i� ܪ��[��xe���	oW�W��s��x�EF�P���f�	�G�q� ���a�{��&�kc������=���XF��B�>�i�e��?�$?5�S���ތP՞���v��]dN�_l'�^p��c�=Z��\�+�;�6�'A b[Ĵ�,%��3e��+��&����)��؅Y� l���i�>�*#t�@>`�,�ʏs��s����֖�ɍ7^��١��z�F��~ϧ�M1G�!xY����G�D��RrZ0�p؝��KO�ޟ��h�
�.�*��@,ö1��Դs6;tW<@&,W��deeϑ�O�<���B���3\+���Ԟȁ���PQ�$ơ\�
1����"������������[�w� ��_��m6�:W~pW����� >���$�Q���$÷��ͳ���?�`�b�l�ܥ��3�Nnr�-�pt�옐����>��=
���J(�`�"ں�ܶ��v�^�_d*>����)H)���\�||�>?| ��%W��~t*����B�s��N�.��[$�Nﶟ��F{��B=�60�Q����[h�`n�AR=����@KN��	�o�5	���i�PF����S73���G	h����w�{?�zw�$;��������|^6��~g��O��b�o��NP3.$�>U~�i�ݵ@C_���j�
�,��7��y�pр�6���=�����s.4�N�_�]��2ͷF�I7�x��� ���2�M�vK��L$���u�Y��:`7l2��tMw�@�I��\2��}�+S~��N
���ag��y��r�*���tSs�����| �Z��լ��
$�8Ri����n�Cz�6�]�	��/Qg�+gH�mED ���!�5��Ԛ�LĤ5��
q���EJ���%^��	���m !��#����R.!{t�����5�[����j�@Y��K=c0^v�b_@^�_rmOY2�^��8M���g+kT�r���Dt4s$�6d��ں�T���:g��Rca�t7"��yxxL'_�(;���d>t�؞�!3�$�N����Ǟ�x>;�U��o�u`� ���)�L��ǜ>��D�u�W,X�SK7�Q��^6Z���q�j7�9=�)���� N��kϭ�ў2�@�qժ�I)�PSξd4�<���q<����������F?J��p6�PeM��v.3�D����Et�L�;�D-y��9���wd�)���@�+؟�T�{�|�u���[|+j`�oX�Qc��M�Ҙ!p�=����*ǻ	vN����1��?���G��n�neZ� a=�s�â��ׯ�Q."����&j�խ�VNʒq�t����r{���G���O��BE �[���4��k��T�j���௘O��
�;i�'�g�w)ֶ��k"�z+�}}�v�Tk��=������v(����� ���p���*z��z���K� RaB'�5�N��]�\�yr���S�?��$y&�4��v߂�d�Tn���S	�����c��7p�����7�ꅅ1����C��{xߤY-(S���d���O#��J,I���צ���|mƙ���$�Drܙ��������'r�b���t1s�k}�'���F�񌇋�68��
�������.�J7�xQ8����ܳ�F��1Vy�H�߯;z���w8h�Q&9M6�<�]�F����k,�-\��@�A����fk9� z_u"��a�wW��JH��)7Ag���V?I({�������{c]{�n 4�*�l5zZD������%A����Ĭ����Ҏx[@���$� ~I6_���V���d�������߼�ww�$�}:K��4-Ѐ�{s^K����L5��6gv��\(w||X$�}� � �z�OD��GN�я���j����{�#傋}C$T#
��\��aY���g�d�ͥ�)�1����NOt���4���lڻx��vi1�=��HEx������IԖ��؈��cf�70�Q<\hO9�ٻ�c�+�̳��6��N�Ɩ]��<���f!�1�"��/�aPcDo� �j.����e���D�\U���JD����E�\`yH9�L��KA?�NO��C˳��=�u7����ڻa�'��a���m�vª -_���C�\��p�l��}=��g���f���4K�����X2;&�Ű>��6�;�ձ��r�-���{�dP��v�b��SN����ꗟ���Y~�<��9"�0�\���>\���w��;[����S(��fw�r��Y<�,�PUJ~� dS��5�1��G��~|愞��>���o�io`8E�L��;�'�k~�w�=���D(q��K�6?B�׿�Zn��L֦����H�v�U���~���!��;��MB�����L�Н����_����IX�e��e�EuSk�W5�X�s$zt�J�Cl͊���4�e1�?�*���:�+����,�P�a��Y�؀���F���oT<�[�ne_s\���/�,��K�җ����Ir�i�}���^�����O �i�.(Oz�1!�g��>;�o�(-d�l�c����#�A�Q#�����ZO�*�	A�$R��]��l=��&)Ӄ?�4��2/}J���{� ����a��ۼ����i�%D��@�,�t��V#�(a����F�%Եf�)�l
�ߺ��@%{";���N  ��h����(\�
� X�]�ͯ��a�陰��&�!�2�D��x�k�9�5x�^<p�_�]c}f�<�P?�t��a�M���W���o�9�t>�-s��\ S�sw�~YD�	�g�B����)Zm�b�@�2&�X���)�i��w�P���<7�G��̚�۹����7S�k�ͯI
�@d�B���9V�Ց��q�e���2%1VY���c�M��1ͷǚ�7�v�c�+Y(�27�/�����!tA��o��l��짲����'�ާS�lz���X�g�(�=Q�;Q$%�w�e=�i��C��
3�jF�~��0VZm��.�)����ذ�5�ʮ$��,��V��0��JeX�"�u�!-�cV��M��:�����CgV,��ge>�<��i��ߠ=�BG���&��ty��f�xG����̐����I,X��㪛j������H��'��ǥ�>n (�0c(��f���9r�����7Dܖ]�$<-T�q�.D�rT
��opE�l)�(p���m���OW�޹��5��u�<��b��, �����G'ʏ����	:(��<�#�؅�<�	�:�?z�m�>�H���-{�E���e��t�ڟj6Dt�O�\<%�:�������{��������k˳��c�X�vln[`u�6&�Fb�HAI��Xl�ae��s�;����^�h��o������g
o��x��f���АJ�{�%�_����� �?�`ػ�$�[RI`k2֦M���`���gxO��
Z�ez迋����
)-��c���V� �_�g��rœt����hrU��3�pM��徘�~~�U!2*�Aj���H�7>|Si�|Ǹgc�0HI���!�}���OT���Ӳ�t��k:�t*��S�U��ƫr_į_ˮnr������F����n�r��Y�}/|�υtGM(]�?�[���R��SO<j(%b#,�@t!xR�-���Y��'!�7�	�����e���,'��A>yش���6Gb�&)�����{��7wí��[�-�tm����'��j��mU)��e�U�1߸.�"� K��C�z�[����s�'�l��;���}3�)�v�"��,:���Y-j��7@��k�����z�!| իL�KE����,�;�\ɵ@fD� t���VhS��=��i?}}r���:����Dc���%�'�Ye�s%)|K˵�y�iِ��	)'y`��V(Ab����
�"In6vp��,��eRe)�-�I}��'aJ�߿����?�!Ȳ��mS�'�'����~��ڕ"��)�u���yI��q�*fa#wC;e��w�V^NW�.�ɩ
Q;���
k��I'�W��
W���7��D�1��H�Ԍ-^�^l*�>d�*���{JU�@��ڒ����@0%$�İݣ7���ӭf6�����ί逪pt���8��:�-���՟��,�Kܳ�o�sJ{���x��5��GL��h�W*mF)�P r'>G�<�<b�3���v�(�5Ta8��;D�@��6�u�/$�Ig����|��e8�qh�i��Z�M�R4�ip� u�tak�;��Z�i��a�UwFk�&X�b7���I"�Eg�Dq��?}���C�a$�CfeS���v�ҽ��R��w4���������ml�Z�����[�A}�cɝG0����X���_)d������&�(��/�&I���u���<���^ڢ�{7���ZsA�l�]0%���h�8�s�P��X'�m�^�-����Wў�Ȇ͹�B-��A��1;6g��@��%l�d�׀z�@��fX�x��vl�K���,O"r'j�H�����<�~5��pl��S +ſ����w�V���4[ �fe�Ti�}tC1D9���)G������;�e��E�����l�{���L��Ћ��|��50��X�u��]I��K���b�\���_��
�7z��n��;�j,R�����<&C_OA[�I<��A��"MnC��0_�⤻�و�ޮAZ=��$%�N����19���ؓ	�ՋwW1�����UH�V�I��m��r\X_uI(��?����+)��*�d�壙�$!.zNذ����N=�ǫh�V��ϷR�������k@���!�jG��K* ���u�߾�$AX��K����f��ϔq�B/�p�ёE������WdK������	^`-8:���xl��K����*��ɔ'8�:!�������7�!_�v���v�'=���F���<w-;F�p.Et����[�����L-�%�''���7Ypv/�'VU6&���wR�!�)M�7��Y/��r��Z�V�\�_�~��?��q�?���(s�sn`|�$��6U�JX�z�H"7e�_�б��5�e��Ӛ�D��;	����]s���G���!�a�P�������f߂%�j|6�j�^p��%��R5�S�b����h9�j}����Ȑ����p��(g�Ō���̼�ю�g���E�ƶ���<�&͆���һq`4q�Mf��,yBt�a��+m�ڶ@�cў�i�iX�h�$�v�3G?���<A����e���'�Z�Z����F�ō��g��`f�s?
��]�� |�6��x�]��a�ҟ�����}���z����I=ˬ �չa��Y��D��*t'L�?>�棎���=I���	N_\~ݘ����v4�eSoHqDZ���y�z���PDU���5t{��>H�\*1����z�	�*"_�����L�!�����>��~��eô�pȦn\�֎)������,5�R����}�>��kI��kt�BV�ɫ9���1�;���@gvh@\�=��(��~��I���rOOʿ�����կ���߿��]�6����C��mY����������5�d&�X1ӄ�'����⥵����ݏϤ�[HNu��ѫu�!�����M�*���"�Fv&��������8><�/5�-l�[�m�x��c���!�g=0  (�*<��X�0`�(%�����(��r��w�xq����|�v�<o�J{�;�A:�/�ܧX�����Tf�1�����U-�� ɛ'ɋ4ck��q���������,�L���Uz�u�PVN�k�<���/+:D��ߦc�Ñ��Z��lO�4�`w++(�rzY@@ to��
Ao�<��%����>
إi�3WK�'�O`���I'���5�a�n��̥�I���7�ă���ݝM���i��+����SЩ�9��ϰS1֥�_����3Ks�*,��e��h�Kk�6'88�� �e�`���NVz�=f��������G����<���?u5�	���,,T�;�N���{U�R67�����6��A )�E��ޘ?�J$E�nZ?)C�e��8�&3�U��E
/��Kr��K��S�U�Kz3�Gi��o������&�/E8<=�b��:8O崹q�UW��`�o���}q�'ؙ+3�����M���ރ��߸ͭ��S�S���~��u.��.�R��k��H�)�륚��G��T��lݘn��[��<��l��+�*��3���=ϸ���g�O�GVH�6�9���C���`���?�p��x�rJh�|���S�h�aW~��.X�)4!���7���1�=�7��c�mG+xe�lڍ��伴gnE�K)�[��rV+�#x���T�\��'m��ڜ<ɕ���ѱ��X��Pӭ��Ŕ{9��H-+����5�m�ޖ��/}�Qqϒ9ޚU_���t̃WOZ���$C�g�_����ض�)�X+��(~� ʃ���)P�?r�$��_�$�|b}�-�Q� �nҀ��`[�nҚ5Β*�`sz6��`{w��{�e�|�(� 2Ra�V�^~0�3�xkM"|���g�,jH�`K�#��g�,�%�=���#���_�&>�A��O��RS&�N�1]�h�6]�zٱ��v�{��D�f1��ef���ᚚ��܂f�F8�>�6���cp ^p*��0jedݖɋ�y=~*��:E��'!#R��}�YҾK}�x}9W��,��'�S�q,�������wwvpڪj��.��~~�M+���*�V��J�����X����1�_�Jg��#�P�S�D"NPWBϸ{��&I9'}N�Z�_��DN�����=۹75�E��X�E	�ã��o��M��/	w+���Oz8��X��'nw_�,?T4����@ҳ��%^`��@���-������V�����#eecf}���l�9��t��T����x��	�Ϥty��$77��F�[����Ҷ�2����[�⇗:�~o6N���$.]ힱ�t��&� ��v�񙛝��M�!9���AU��Wh(�~U:`�)w?���A����K(�"����F�+�	;�9ztfV�k� ���֚9"}�	=NRH�����V'�C'���)�����r!��{\�d�t]��g�|Ɖ�,���sU��j|������M�)N�\S�hXKW$���C�(ljk=��u�I7vxl��@���qi�<��%�������2U"
���03�A*��'�r)y��n�yV$g�0��gF�&��)*vmo�4�(N�����D4�i6F�=��|)�ȷ=�̄��]nأ��T��y4�o������o��g������56LY��z�3��'��\>p�"e���������yR����u�H�ǲ�P�1�����`�Y���o�|X��I.�,�5��O����/s��P\0�F(��D��^dqdw�,&D�z�`��C��� �h���q��~m��hO�BS��C���]g����,�45$���jғ&/E��s<}^M|	^�l�RZ�5ڭ�;Bw�$��	�޿�(�X���iNi��,�D��TN�!��8�#p�]�Ǫ�'�J�.t�&��]� 4:ofB<@���rȪ�����ϖ���6��A�Ӭ��0��Y�#q#���K�����x�s���w��~cc���@�+ �N[�vͦ���.u�9�ۘ{Hm��xH���(��v!�I<��!�"ծyRS��
2Ƚ���.@+�䂍@�d_d�P��t��
�M��-���Hq��Sخ�5f��@�Z<ՏWK�+G:k�ع���f�^�%va�J���$��9�Wᣱc��J��
a�p�)��/H�M�΢��|���X�X R�����՞ڗ6���Z`�G`�%���� 﫥D�OF�þ��k�}C�Pg휳}���w�<��� �RϾB~���J�pF�lM�z��w�^���9y7�u�D~g�J$S�EH&;�z�K}�6p�k&UD��Kb[c,t�/�~6�
��3�_�w���<">��0�[}���x���N�E��b/�����$ih��O��>���ϖ�����u�ik�%��߬nm�8�������p��NL�݈ryY��p�	�`-��{��HQ�C���y@Cx@n<���<�	ߗ|�@:/�D>�M+��C7����#����qH��A�3���z�>�����SV�����_��M�|�gr�Y8�iD�f<��p���@�D��ט�\e������썴]UX��|d�-D�p%b"X����k��D�������Rɪ���t�N}�����u�������V�x��u�n]5�|Yp�VF�8�܏'L��F������i�<>>�}-3���<��&��歧kN�Jwױ�2f�GSC�xJ��� �K�
���|M�lT>r���]�>�S�ߊO�J����w\A2c"�`��	�R3R}���f���`��UY���+��("N�W)��?_�*��
VK��֤
�5��[��\R;u��%=�q����ɹ2]Պ�q�F?Deܻ���מ.��ollB���w��G-^>Eʰ�8����H��t��{s$^������v�*���r��F��o�E�6��b;���$sڷ�sD��cߟ�bV�	��~_[�?��;'���ˑ�?��#ۥH��i}�[�`!���g�B	;r�TsF����`/'dff�~�IN�o�C9�ݱ�l��[-W0�WhO9ŕ)��_%�zqmm��t�y�n�R+x���#-8��u�N�V���D>qS8U�˒0�2�ɥѵ��4�/��[�l���NIc��$d�V������im!UUݕ�N��m��7��^H�]8����[U&�k�`�3���I�Pơ�0-���L2�nVœ�b��Α�O#�
(�nƶ*7m�#�O .���8݅�(��ڎ�VJ���U	����`kF�؃;oi bV�ɘ��{��+p�z_���"f��fi��h��\����yQq:�/uU���p���.Q�D���LW��J����,��_��U��E|$*��
���&��v�� l_��݄�FI	���v	��m�gW�8�� 5�q)�B�����bDMG�S���e`��t���ڍA�|3���������G�y�|��\.w��*ɮ~N��w���R}��}��A�W���\^������@��*�η �a8�������m(�\�;�d�nǑ�vaF�R�n�O�Z����h�M&d7C����ɓ��~aa�YY�i��p:.�3�S�D
q���6P��s�K��S���_�E+�Z����`e�/�/����!�yQ5��5�T\�A�撩4*��>%zIY�SUJO�����������%%%�R��t����T�M����"s��O>G�������."�t#]���HJ����K����(JJ	K/�t
H��.%)�t/���������Ν��<�ܹ���m��+ݜ�U*��ӤU�4��>/!d7���,s=������N=����D��s���%C��͏��P�CS��F��$!pw��N芧r���[+��������Y�v����D��[9����\�A�dmmWe����>����|��s��y�'��<�tg�y���N]��;ő'A��#��њ	�� �N�w�(%���(���TJ^S�����m��$ţ�ǔ��U#i���+�<{cs��r� żK� ��@�C����#V��E��i�F_�|���h�vF�}f�m/��L�~���%����<_��ff��g��9oծ������(� ���2���D`�CP	UR�)����kǴ���f�<� .�K���(3$nB#4 ��?9Ҕ �Y�<3^X_YK͓>�"A
��9x��M+ �%'�Ɉ��=k���ѐ��8G�6��q���m(Y�o
�a�� ����62:�M��xՆ�t{hӝ<"~�g�m��%��fXy
q�X�����lz��O�?��!�x)7h+�u*c:6�����SuU�'�#���;R�o���A�G� ��?t��H��6H9��ʳ�Wҭna����<�?��7J(.�կ�o���J :5~��?�Imy�˹q���.*!�Q$�������U�"la�;����a�u����͆RI����}5933��'��X����zza�W��-#M~���60d����2a�ZfO��5��W�?eWQ�dP��~�Ϩ���;9 I���QOn�H�G���w��z3�=���)������u2���'hUm���v;�-ak�����ηtg��aDћ��Br���k)��̵Y+Ƽ��,f���<u�$�'�,g� ��_t�اII#�]�xj���]��ah�t��A�%W�I�,�4 e�rU�Ҳr҅�V{O (Y8x��YrETP�3��2���q-�,|���W�`}ǧOҽܸ^
��D�ԩ�O��)&2�D|�p���?m�����⽹P��ĽO�=�8jc�?�
}��ocE:ٹ���G�ăc��ui;�ރ�#�k���Ԩ>�Շ��d��&�#�v�ф���|S{3�0��_�i����qEk���8�7=�$�ɕ� ��~�lb��q���$���ؘ�bE�B�Gd$2A��t�vw��*B�æWUQ;=��QaeWi�r��f��*�-P�C�v ��ƾ���6+y�=�b�hSr�-��T_q�_��squ����Q/d���A���K:ܮ Gr�N�7���X���]�{����6v�� ���v:���0��+S7�J��1�ʻ>Z��FrK�*z�|��8����_'ߗ5�w�"kt�aMlC��O��d��mxi>L��&B��Њ��?Z��C��=�� v�߻ᡷ-�~y�f�X�:k.^Iى���sI�G]�n���XG)�Zz��'���;NN�aE�'���}@x�D����"9(��(qp� D����4E�|K���bW������|�0.k.�Y~��^B�H��~�<�¨|�(H���ɣ��7�/��Ytէ*s̟�O��xƺ��+=�`33�A�י��|��6w��!�H��d}X%bz�]ߠ)9+aO�&]�
Ĉ��+�%^�����r��gB��&S
?l���S<~���[�^�?�@�d�|TPƜ�����4| ��*�!�s좭&D�U�����e	f�w
ǥ΍h.��4ުCުH�}%�妡R'���^z���.��	�_�I����D�z#���r�E7�W���{�)�\ �����3��R#9Vq���d`��B��|@�d�����AP߿�v?���IU�7Ӣ�h+��������3�Sv�F(w��y�f
��eh�kF�;��{��J�,_ҹ����%� ��&hfN)9������2E紧�*�ԃ��KJ����������HK���E9���O+�:i�wF	,M��$@P�f u�L��Z
;s����7�(�d�Y��y��a+�4�b����_��	P�a��~maى���Uf�=RaQK����U;GY�d����w��uH@ǉ�v�]��CY�T��-��4|�K�x��^1���۵�=�����WM�$��.M'(��I�U�����yyv�@��=�<M/�aPnq}�3�����Ig�}��ϟ�6���ĵ��{����;��J�����	��q,Z���+
3���h��i�ӺP�=��gl�*i��8x8Ƕ �����z&����H���Ŷ��b��TBDz��a�L����Ǚ
���k��x>�\�z.<������F[�,��Ǝ������b�YCw�V���c�������t��jE:�L�y�\U�?*r
x$Ɵz:%1c��:g?��>����=-�'���$tD��E��I�GO�$<��� �����p�2�"�Pܶ�X����p��/��m�_�����{�a2����Ј��?i��,�P���]�^`���ͫkj��-l%YDBL�k�YN����O���Ɏ����:dV�1��'C�#嘉M*�:�xc�Fۘ���04�2�"�M�iRۗ��'�]��|\ҟ�di�7�Ѹ��jt)�O���̢K�A��5�0��qҰ�Sp~k���/�<q���?���"bg���u�P�yWq��s!������o=&;�]`��J UB���^�O 6����Ğ���Eu����}����U��|������L+MM�i������ע�F��̃�[g���ʗ=�ҘWnKz@����s�RvK崽�'=�h�h7�~��������������qE`V���+�O!AS����A��q�".�����_r��<=�c0drSS��\T�F}'�-4�2�n�;�S�$��N7__Q�l�{����>���˦��*��]H����|�z��L�~Dr��X��̚8PB#�ý�s�A���0�|��+D� �L�3A�5���g��5�}aa�k� ����,/N���NY��J��+)V��6�!�;^��7�L�pXe��E�ǲtX��q�t|o�~�jH�V��"S���M�#R�C������v�V_����!�5���i"�$�瑀ω�1~�l��U�~�qC����B��x?%��٤	4�z����+׻/V�W.�S����g��{k�@J��ʠdg���ɐ��J;��pq�����|���m�т>@zk��e.ψrB˳ ��^V��	��� w�5yrR^(���	�����.���q,��������zl�̽�TE*47�|q��N|Ez��y����m)��e�k�X����R�>�91
�i[���ߜHqw0,�֧�|:����ߟ�<���B]���7�jb��S�I��-���R�8�k%O�;�6�=*�$y,IIh�4
� 8�*��K��r:3��(y��(�LF�F�����S����f�`�_�f�6�]���0�(��0(�??���a6�28��b}1��"��c�X�"�Ƣ9�x����V����n1]f��ͅ�Q1���7U��9�?�f]I��!^�E��^���D��e �����\�2^���	�	~@T��.�4��v�3I0Q�7�ka����0n�����9y��������q�ύr�B���+�Y仓�(F>+����zXbzdjj�	��L�*	����!X�G�/# w�K嗦H�����=@������:׿�V��l3T�e&��8J��:M����]}�I�Q�ۚ.Rbv�P�"_a��[z�lk	�i��|�$�%�R�{����[���Ӌ0�N�v�0�Q+�U#��l�*66v�ތ�V��fo��o'�]@���W9�K�R�����T��hN����>͡���U�w:��2�S���2�� =���Gl����R8�Ks�9����a��EQ��'�z��nP�7���]����+���e��~J����~��	+��@X*���b��̌j�#P��[��)rξY��L�˒py{�C����U�i)����5LZ�ꬋ��`^����M�=C�����ќS����2�/p�,�]�8��s>���i�k �2c�@R�oR��#s�����U�E�S�{�o�]�1c���
H�_��+�<��/�v�N#A��a�	��'���Rv��1�A��'�޺���]N�ԙ��U�t]|��� �NL�Tץ����������{�LE�j~��`F��7WL�	:Ó�X$����"[ת�k%)4�P���P9T���@��a4��OV��vi�Lu|;����t �?��պ��*c�d����~��܈���i= ����0A8�{�+ŻK���baqr0SA	�E�>O�?�:����%���o��_��) ��97U�D�T��!�������S.����W!�,,AA-���a��ʡ���-�s�����L�y�~	����5jS
��N�od��kMh�</�I��*Kj�Fk(�=�׫_2s~�|$�'��!�euZ����D@�=���;�� ?v���~Dnf���i9cy[ Y��239r�f�zv/��[�1��݁_�E��e��8
�
��K�7� �ER%q�"��}���Jo�nE�*�n����P���o$[�/�s�붖Fz��5�҂���r%kٔ���^U���h��v�$���{�/8��yl����KD��E&x�0c�بa���T64��W�P����8�L���A�ǫ����O!c6�O8 =���KO�Q�~��VwT��kw�;�m��	�N0c�z�Q>3E�p=@�u�#�f�}[ΰ������I�N���c@�)i%9��rty^�4��K@���V)��cwW��~��+ϻ��~�кO`��i����c�Ba5�O�"�����z绋��N���6B����jT�fNg8�W��[�k�A�W�߃C��8��"���c�l��F7{�X��I(�3�x����]Z���Y�Ã;L��2�@P
�5;�HM<�����x7�;y�9�c)��j�
�X?WQ86t.��\�~�~ �e Iw�P/zIpx�w�D������2������ȼZ3�#�+Dj�-���Q�D���ŭ�`_8�ց�%w_��'�>�`I���""Z��YP�e��췾'�=�ߣ�{�����07�yF�K�9������	E�Ng�Ӻ���^R���B�tk����7���Ӗ?5�7b<6�!���)Х��fu-gV���!�3�1�}�D9��PX�V'C&4@�O�V�D=
�r���a�S�a�X�V�$�ٜ��|�Za&�MJ��잼�~�?��M�\�~V��''i6�ٍ֭��Z�4���D����I�
�K�S0�S�S�%��Yxy�V�"+5�����&�I׻��쾂LjOAb})�y��q��>��C�Ahs_ޤR���}'�u��t�n�����@�7~$_��G��NF%��;�T}3_AW=�6��OW�L����z����R��}[����P��G}��'�޳W�y\s:��I�IO;7��4}'��᳾�7|�W؆�VR�e{1��Jw&�9W@#C���H��G� ����tjJ����c�֔��Ov�p���fn����T�=9����Z��R�`\/��y\�wH}�j?���U�N��%�@�y)���C6����w�T�\#+J�m�ɽ�K
4�������
�N��~�b'�ؿ3��M:� k=�Fퟔ2�[��J8�U`��k��o[]����Qv�z��vmhh��z��_�)Qh�: �����!IlL����߇�o��J��_1L8
��J��ޫL�̣�p�bX�s|a��Tq��AՎ���{��l,���ߧ��zi�W��''�PC���C����
ܭ��x!���o��s׳���?H�7{p;KCތ�RU�iKL�N�yw&!3h�d��%^MC� �?{#�֣L�y��t\����I�ҵ4�>�pQH���H���9�|�N� u�V#��Z�R~pdW�l���E'���������?�����F�=���hV-��I�X{�Ի�67��D�b�cV�\3&�+��~����>�ݙm-��q�]����a�I��x�576R����]~�/����CH��x2�~3 �	
��rv�e��|#U~���,��H��r|�>�@�#������++*,n�TG1��n�77�������
�ٖP\\�u��HK�,����Z'346�K��{P�T�C�N��;/.���3��Z׊���s�-�M�훭��r� �!�rd�0�ef��I\��]pӒ�b �n��#ŒGY���fN3S䍶�|��\�[{���c����
�~=O�������+N>��\,xdu��Z�Q�R��4���~��� �O9H6�+��?['i�3��Q"&Ǥ���z3H�cI	/�����3,�B�E��FH���tI�޶d���,A3S��.�T�/�e���x���UQ�ˉ�ç����ퟥ�9�~O�� �PYWgW������G���K�����o�������nN��}�1���Yh0�z�5�r^"x�9xy)�U:��S�uo!��S���C 姫'N�6N����Y��@uuV:�uR~(������X�����H&Y�_U�����o��"I�S��u�������4>�U�4ޔOv�N����9��1��[__oPs�tJ����m�t5(8�X$�g��9&>9'��K�!d^/��2��05��xX.���s9[������9��z����W�K��qo��c?��=���N8�������`�\ӁM�����rv���]���U�{ɪ���eѩ�0�A���E݌ȣ3�!�s��5o�W��-�P�^�1ˆW��� �wSk��h �h33���,my)�jSUE�cnBf�%aJϺX�����?>[�-6��y�j��q�$%5u���up��"��
d2��u*��1\�,��I��v�X���4�N���J��L��,L\:���t�O��m��-�_����,	;���R��F�u����kà(���iW��v���]����5܂Q�{;54�8\O��fw� \�U���듛��K���e�����_�������egd���p��*���,��I~_��y���ȸx�B�_`���}|0�0�l�F���<t� _�� ߢ��ak���!��n��u���S�g����LO��]W<ovM�H���W���x)gn�U]]m��Է��i�e�\�>�A��F��O��=�h�?Z-8|�}Ju����Vl.���V�C����.w1���5�>�;LF~�)i�_F�sٛ�3=}�r_:Y�Ԇ���who�>0���\Lpq��y��q��{�b	6�7� ]9���q���	*�~���+!�ĻS�j�Rm��ǘ�"��Y�D��r_�+P��X޸�?0_avј 4�0��������wB�>�݋���ܤ�̵����R�w%�픈�봪pH�;P"J����k~�Yq�M�f�h���"�i�JM�V�e$Hօ5Id��#@�]Igu�)@�n$:Z����㐬0ˁ��Q]�̂����U~��-َ�$J떿.VVO��7�1<j0��~�����-��Vr6�!�a�S��i/�~�5c�4f�/al,���"��⽼�	���j:�j�kT3���M�Mr*��<؊}f1��<$�U�~���jໍ��+s��8b��aW�E�V�6�6��u�R�=?2�x��M����C
�Emu�ѧ_���=%��3.ӯl�Y�l��B��4�ÄOH�Ŭ�u��[Qxs�*�XF�����I,<������,7ifO��T1�=N��F\�s�Ie��-,�����^�qz�	��䋪oP`��OSÑ�3�F�����&�dP��](KF�(���m�cg`ȹd8�v|�`:�7������q���^n�D���@rK!��>�8Y�ڥ8���7��q6r���Z��w9�������z~D"�h^ب�uʎ��ˍ�F}�_T���%3W5��>�q�Lv��
��7� �����ͺ�(��،���#QO)�!_��Fo��/ˮpN���z�Y�F��9d�_�����ir5�"�L*�}�!����bɨq�*WV�s���?0�]�N>2� s
�2�S�6�mM]��ߚ�:3s�'��	lD��S&v����Zf�P=���1�ۡ0�+u�ό�����r�;�˙t�ΣA�3#^Ϗ��OF����
����~
�N���I��D���`�?��	&p�H~	���}A���q�[�b��:y�.U�6���'
x���ׅ�~,��2+�h�@����XV�
�����y�% (}wqʁ����,IU�QH&��UDЯ��웤��Mp����(��X���o��(]]wث����⫊��(�R���G��>��a���i
��b�����o��2�Scs3��%>���<FBL�$�}�<6�ۛ)�����_+�$��h�JL�+mD5���w?Cw�lW.�F4mL}Q�?�~�8�>E9�G��6���(	9?cH|>��M�v�@�MAِSKuI��މ���c� A�T6��	���<weSv�/���Փ'�� �^��4��mZ��5#-�h�tP�-��o�ow`����ԄW�ⷢ߮z�W[��tX��$����vǫV��MLlz���n�F���V���R������Jl���h�d���[v�/u��o�i�]zV��K�@�̄	H�~�NX#cEA�ew~ff��kYk_`q��R�/�|�-<,��/P�EAi�Sp/�7uE�50�T9��M/�M5j!��R����bfH�Qc��pH��i(7e�!�� &S��˨hu��:B�qH[�0M�BYO��R��m�ST1�ԯ��HI�޸�ΐ+A'��O��	J\)�����`:���a�H�Ϋ���{�v���1'����s��a�8/nK,�{=/@��`�4f!����c��M�Y�"D�n�<vs�?8�?Ľ��� X�DM3�مE�39ʒA�_�vM���AU)_j�OX� nIE?�*'���������)ۈ�����y�ۍ��Fl��0-)z�cM��?�L����6q~A	K���W$'�A��T�լ;a6�N�s�[tV����xL���4��E�!��Sl<1��gݨ3��k���а��03z�q�D�̅��7��ք8}0�&:\�Y�eF,S:~������x&QrV7�.��zq�����ܬ(�eA>�"��#͐>�T#�i�HB5u#4�,�n�V�u�6�:�����/p���z�t!4#rG_����!�ɂ�~��z-�u��"� ~�a���r�/�Y�؀p�WElU:K��NھbR R�C,M���6`���<ڝ���j4D9�xjM���y��t�8�+!�l�m��5?�[�|�K��:�}����vzJ�����"fØ�F
��ϽI~ҳ)���y��b���3��0{�Y�WލT%�^�~%���m�����3{��H?�½� M�uN�!<Is�#7��JE! �(1�#奓@|�UݏN���k�'!�]�c�_��DQ<��<S[�|���d��Ӆz�j��J�C��$3Q��r�=���}�w_�EQ�}Ѡa��#��ݯ%//I0{�oH�����q
�v�:�?�t�"`����
௼��F�c9O���/���܃v0�h��x� ���j�]y34 �ϥ�α{	\V���SH�;!>#�,�N�|f�`Ԇ���8���^Պ��/�Y h�v��j+_T@��W)�
GuاoiL�?VCRA����G8x5�ix���M5��l���sNz���
~����>WN�-s.*f\vK���Ɠ�u���%%���b`+�o�- ��]HS�`d~��W����T���D��)el�h�gz��׽癛�?4�M:z{f����4�F���	}}�'�06��v�|��ڍ���z�N���F��^��*�a�mt&�S<�V 12��<�S�/�
}`��AF�8�35=@��b��P�H���
��O�dh"9A� ��hz���^�pE�#=P7I�٭�Yn9g��E	M�7�D���?��4��V-\�}�dH���_�=�
��l/A��|1�/����Î�i&P'�/�t�^��]:fw��^~�b:;���k����9�k�/�� �����^0tZ^����� "�#��i{�[��;���]J6J��O�(E�E���L�͏��Z5}���R�
Oo����l��p���i[y���I�c`�;��Q=$ƥN����ԛBPqbCK温�ow�H=@�zn�ޮ֨#�hs��@jx&IB&=�3�a�����}�X�*��ԭ�QRRo��C�t0���~�l%D���!9f�9�Z�3��a��w��2�nÈs?��)sw�:;-�Ћʉ�����y��v-��O����^����Qra��hhX��׳)���=r2��3V9�~��Ǟk�& �u!N���פ����I�MB��Lx�Wg����Y^��m�z|=G����n���(*��x����M 5��k��� _N�
���u���A��!PX��q� [���b�'٣��a��T9s��׍��9no:H��c'Γ�RFْ�l�����}���Ix��,������%a��ӯ�E;�hZ"���r��8ā`�I�tjv�����mI��
㲷>9�^V�]��SoY�.b.��Yj���l��>p0�>󇉀�)2���(��ӻ���^k�鱃Mj���d��� ���2���?�Ӷ�����Vr�{�C���;q�����g�9�;�_#�g�+KR�[�W�?�Y�����6"�$�Bd�Z�*�Ӭ~��@mo
��؄�֊��X���b���_����Y`B<�ă��FW�j����ꄸ1�)��̸kޱ��V��������h�}b�i,�5<O`�t{���ʐ당|�ԉ���)�i�\Y�Y�����]y����{���(�&�S��9���va��ڝ��x��	KKr���2�=�K�>�v���2T'��� 4G���T?�F��)�zq�M���VE��$�e�
F�_e�rUmi>��~o�pѩ2�$���A-�qߔ]Y)`a�/��L��'>��K�E��Ta�O��P��E!�2��'"y!@���L_��'���y(���'}����;9����؟�/;=���͵�e������8�B�`t�R
�wM�Z?[�U�v��W(�����F�W����@i��!��ay�[�����0=W��q�e\J���d�ȸ�a���WAo�q���G{g��R\c[�M^�>��@o�<�I<1^�`�ɺE:��n�����H�+��cE��֌w�ý��-Wq����V���{%3o�_�P+ao�����ݴQ1?r5$vss}~6�I������bo�z�G����q���_șJWJ�3����ย�GDj��BmS���+@�Q9l�KQ/"ԍ�.�ՙU8���b�5D� ^�"��w�1,���[{5��?VkC�n�Ţ�#��O���7������F�C���}U�҂�E1QM̽ny���C�l���O���%]�8�|��JW�ٹp��E�7������=���.^���my��=N��UQ�B�lTߖ��KcR�Xw�p1ԣ�A��.Ja����pzo#��i�&K��`d ���媟l�gGϭz`F��-�vwZ��b�_�'��k���5��'�fsw�2
�`-�w@��e�ט�$� ��͇��ݷ*J�Q4��l/܀�5ݛ�U�>�����z���t�������(��?�u�;"e	��qj���7(vS)�.��ʶ��:u�9�A%5S�P�bQo���ׁ������D`I�EupK�6���2���4�Jg[�l���*�Q�$������Z�ZiB*�r�91�iq7b�u0<�<�f2u�"uڱ�G;c0J�)hv�MGǙ�x(u�k�o�"mo�b{���n�!��L�gV�]��{A����(�~��p�K�}����S'�*B��4l���>G��.Ԇ�˷�k�E�t���m?m���E5?�S�e��S�[��_]	}y}�e_�jPgG�;����ț9�e]�N�3�'XI��@��Z��(U��Z37���SP6�DJ�8�\V��"=�$!D�CNL0.k��cO��툐?X�ϬCsJ�a���/#�E��݄l�l��vq��򉱘-zl;�LŪM�M�6׻��J�ڂ#��7��>�	V�p��-u��.�J O;p��k����ٛfx-�2o`s���n ^��ڹZ�ǯӀ�^eҕc��73����ڷ�J��r��2ɟ�|�J��?˙�Dg%��KWא���f��dG��3w:��*j,��r2i�E����]P�m�L���$�)KP&f���
@F�^��6CR���L�b�u��l�&|ѱ�V�� x{
"9D^��fG"d=�?�"w�a�&�G�%����Z��.]��mp���O^��=��Q �8��<�uN�؀}�2 l�+f#�m�:�ރ����J��3�2?IY��M�
���ne�/e�!˾ŝ�.84@aw� ������PVM����kO��^�/<d�N�5s�9N����e��O4�Dʹ���C�&�[y�D�@�[�(U3d�	)- ���wgb�A"����Л�o%�����>"������C5��]�N��b���ŇL����:(r�����%+j�,����SH-��_q�g����G�����m\�ƒ�H�tV:�5E���CP��X��c}��ƺQ�UyiA��an�ū#��+��R����u]* �{�: ��3cv2����bTء/�&�<�"�/eP#é	��+��UM2 �a�&�5�vb@�p�]�dB��MZ�)P��������2(��8���'E���T!['���f�ɪ'@I�X8`�{���@�t��A���[ǣ���o�9�	���f����X5�9�/f,/����]����f�J��Q|c ~��۰#< 6�pF�ӂۡ�I&r���ȇo�zxx�DL�Ɓ����*n�@�d/� (��5$��q�b��S����̤s�#�䝁�,��u�K��MB���-g����r�M���6�ۓM�p����7�S�hܦ��i�����g�1iN�fH���~�/�����LlaQ��L�.b n��B��i�UZ�0�i�_��~�V$�q��H]������EIxD\VXԣ����OJ���ǃu���dE"|�?wށ��[ZϢoR�����ֳs�i�7t7�	�-o48%�u����n�YH"�k�Gks7�6�~�)�� �jR���/�FP��ԓ�,��I���c��csĩߎ,}lo�yys�4s����4z��\tw��l>��6���+s{����$����A���!��ɱ���ܤ���9��zUX3�q�.�����_���n����o���2��S�Z-�L��,�%w�:+���O��S��BXi�;�����d2�P���t��X�R4��L�Q�/dL*�.[+�د׉k����n���g��&\ ��Z��-f,Mcv*��u9�l,ǩ"a �x���,��o���Lihii�|}�
�T�C��+U��RC�6d[���\GK� ����1+�f,wsiqY�[����	& �+l�
<�"-��9.b[m��[\��^m��lP�5v�$��;��'������U���M�����	-gK�W?U}�7��Z����BSO�Oa~�^���_�%�W
�[/���w
@���A�;l������>����6�y���S2�Ѽ5�Uv���ԓV���bh]7.Э3Ίy�?7�'��c��O��K:L�7;���,���� ( G��bo<����u~Ŀ�;����Ŋq{e�͙Ok~��avO�BK��yuKy���IɎu�s���A��Ϫ�G(��vC�f��#��a��L�^'�\p]	q�yk�����rצ��W=��s$W�jM�Rsӆ/��q�W����_�g���Gm��Ϗ�Zm�r3Œ�O�g������@���E�e� ����C�T5AT�"��@j�;�rx�qY� [�L��P��+00��u޷���-YdksKNj����,Utu_�>q|� 6��;Ώ�B��|yjFo+��*PR��o���82Nca�%���sF_�G:��#����rc,^��v��r���Q`�s�������]Di�����l��YV^A�#�����[�_-k1�@�{3��������(���;�ަ:}G���A���<ۅ*�N���~�D�+P�1@��o!�o�P�S�!��f��ld`R����ϛc�wv��]�5j����=�����E>r��b�&t֏�9i�[�>3_EQ�7_��46��ޫ��I\��F�Uߜe/����A��7���k�V�����S�Q��DkCC+���9�֫���`��������:����	����� ��5�����ǷA'�}�^�|{6��=�8D����d�,�ۣ��.::�����ͧf��c��v|糭�s�Yǝ��2�jtB�l���1Qr@s�]��'��焪�VA�ˤ��*N��A�r����hu�q�­s���EG6fj�꓏=c���n^CP�8��sٔS�����Y�;or?@k���@eOA��e}�'A��o���	���?����A��M���Q���-�2�m1]�n��Q���w�Z|u������͑�H;K��_��{�-8�J���Л��sް��wD)�!��'yo��Zi���
T�}�&����K2��.�܇����p���эq���������a�K�)un=5�Q}Ae�}p(�)ߘ�zĸ�Ɲ���UY�Y��T�5�C������8k��ě,�B	W_����=�����1^�~�U?�(�c{���7�:�L-~TGw��R��u���I����+#��d�T c6wa�e� A!vD���{@3����At�����ʟ����~�ũ�=ٓ!oU�ۛ�>�@�A��^��~���)u���O[N�8>@�6F��҃jbﵲ�������X����'�N>�X�����0�c���,���wCtV9��7��4j�v �_|Y}-tn����n*������v큸����V1a����G>v}�2bZ�G}�?˿����Ϯ�������0�N+�&Ű��҉*t}V���~�O3�Ker�����'@|=��V�矞��kL={O�Gh��%SdT׵�N>�yB	�0�`�v�����m�T��8�DԚm����S�_887���MU����F�o��!q���Zn�aN�e�@w8��[ҿ�����Y����R¨���vBo�%���yW D�!� �eQ*	�gi�Y��9���l��T��I�>O��EA��)��U����^��7�C����#[ǘ�Ҕ��{e��,`��rL�����t���Y�!"+�ɱ�� ���ڹMQL�B�k^�߁����5)T@`��n�8�'�7hZ�&�J��l����Lwd����r�H�{E⢽7���.�&s��K�;��폤A��=M�� r��H���Jhe^:���s}�A���J��e>M�I��E�P�^��gs���O���qv�`ߝ{��8�^5��z�@�D����nM��R�����z9��^�8�;�+��NǶ�)�2 ��5{Sk��9Tv��sӶ�=��[�B������nW�$��;�x��=�#8�Ы}����@�|�v7AVs̮W���C)�}�ؠ�����#���n����4r��$$�இ���?�k�R���A0/4Ͳ4�6E:� 9�p�fS����_z[母�&�;���R>>�ݱ�'�'j���6�E2���,o���H�Ɵ�O~;F\�_8��3|�8���^�`����ǽ����P�K#6'�r�7����a��а����o(���Rvo�w�02���Ĕ�2}7m�2����i�1b�qT�N�EO��{�gS9_���N�BdM~D�c�E��9��O�F���@|8X��>`j��k��jP�����+���a4n i& �4&�rs�z޳��̱\մ��>�ϱw�������wCYC%�����B��5�-�k�n���0T�ԥ��v ��}���I�߽���NR�M�k
�g�����:���t�X� E���^7'�r�L�f���8�{��wH�Y�q�P��mw߸�C��z[�ȿ�x���/%�Ma�CP���m`T���ז��1�O�A��/!������ 2���q����ivM�t~-%���#���i+�T���\ӿ{�a��kx��lnݐ�c�Q��n��q��ފ�_��b�,�L@B�F<8("�x��P��|,��}���ا���������`�M�IY��,��DN�X��4��E��.����*6sA�x�n�w�B��^��t���	�鬡ʲr�l��C^��*����ܜs;���l|@>���W7b�.�,l.����ZB5�p�z3x�ov���V�jZ��\�Z�<���ޖ�`�O�3�f��A���ֆ�f/�9��j��4��hNLv�$},���-����=��ٜ��k�Ǣ���L�tu�b��ih��ʷ��_���.Ao�%�*[�"Pe�+H��rߺ����U}�!�PO����Z�sV=���q���z��T*�L�Hk�%��hV����~g�.�����Y��L}uT����"�H
()R�A7̠��tw�tJw(J=)�� � �5��м3������`��9w�}�>����}�T2j͡Wf�\X����v2����1v:˥��y��F��\��䢒��#Th�)���a��F���:�������RX֪�$I�y����@���jB������YU�0q&��'%n,�&O�[�qm��YE}�:JUdX��*�|[z��k.�uk�0\�����"�x[���5�0tR#��CW�j�ʭ菊�	��t�'!pMdɭS3'}e�L����a�_~�v���O��ߠI�Y_.��z�i��������f�%���V���pw���:���Ҭ��u,Z�F�Ӹ�|��Y��!���60�L=Z{r(��ߒ�/��67��n=�x�V��4��e�+L��^���7�ݭ���A�o�F$�a�e�|�b�����28����m��>�榬�Qgǿ�Ԉ��Y Z�	�/��H�dE���dG��Չf>�Gc}�\	I�k[�?>�0�c^�R�?�0�%��
Mŝ��F���
;���Z�ɚIW	����]���S[UEw���[�:V{=�A|���f��:H���Ϸeav�XM'����|�3;$E��8j5�t���Q$����l���;-,Oz���(��ߏ+�7yR�_��r��(��=l�ϧ�:c�@ZA9���������b������骛���ֹJ���-�iV�e��k��gk�+�%�oht@��h�S������<�u:�n�q�[�u��߮7o�J���&��W�!�Xٙ��e/��
i�l�Lz��F�W7�y�������
�ឥY���	�_�[�*����5R\�p�f,I�b4�S�C��o��29�b�3�*죪�Ϩ��5n��T��P K]鋫�G/�S�]fb��䡿��gs`��ÏF�5Ė�<F�,�E��mN��� ˽� ��:������v`�]�_��� nR����ǿ ;6���?ΤčVٖ����e{�x\05�1gL�x*��Z�w4��c�m#�96D|hG�:fѲ�k8���mp��#j	D����ԛI�ߡ��EQ�ؘ�i�ո��=��Y���9�moI:�6dI*�ȁ�"O������(���'���Uq��7�/��#s�/�Ф�D�`[!g�肘�*�Ǽ�Y&n�,7�y7���Y��uhh�Ͻ��.������U+��=gF]c%5��|����䣦�ԁ�����x$K�[�6���cZ�Wώ�ל�<-)��|�٪a  +8h����`WD��ݿA��C��[��_�&ؒ�cx@�!���C��5b�/�@kX��Q�*��J}�ﵓ]��f�{���noq�U��;24����U�d��H�E<}���R]�]ޡ3��r]�%�4��^v�����X�Y������9���pr!����rB㫈C`@7�828Z%����y�1���]�2��ܙ��ӧ8��h�����	փOl�O��a��0�������I�g{�p���}	��V1���Cmƶ0�`�u��+�ž���]@MP���;�XO�\~���'�X�n�R����l����' i��^^�#�^�a�ZX"���	f# N��}��*!�X]}|t�"�z�*��f�N��1
]8�����FZ��/� ֨��`@t��A��������b|��HxL	n�S�Vd��e�%%%��t)B���en���/�F��=�4��'�f��A�#|Gw�i��(L|�~r֩}���N�5������槑�9�G�7�F���)>g��O��u[@I�k�7-���x��i�q��x����=�D]4mZE�����C�.�=���4L+�a���9
�6�P���W+�k���BEmDM���X�ؕpx�O��J{S+|LÎ��n���t)e����Yx��s�Rٲ��-���u���G�<T��Gއ�/��[�o�լҍ��1�u�o�2j�d��;�]?��t��k�H+�J'�z���B�0k��u�9��{Ew+3�b��3�m��I^O����@/;�ܶgl�!>�H�磔K��I�A^�(7��jQ�!;�&0���i�a�Z
m�nǅ�Zl��o`�Dg�f������p�z�U�"�O�k��%��Yg&[	b��٪a�����}T���ly'=��2�G�.��z�)�ߑ�1:+`|��tf��B؏m���ڣ#l'��&���l���A�,f"f���#�Uq�[�� \n��4�S�ssM>p��~BG�Py���Y�W~���\D���$����aQ�>�:L��(u.~.�N@������Tzr��<㋕�U{ʕ`ԧ�|?0��t~/��.Ռ:� 	��y�k��Z,��Z��w��D�0N��s)�=iB[.�S���J��1�V�sS�j��׊I��ϛ�!�[6��вz@�����&���7������� n[|���F�����6?��cG<_���Z'���6�(�^ǑD<�j�X�-|3
8����G�^\l"���w����_]���5]�Ȣ�!�c��|�$Jq�>%i��5��%7Eǝ15J��:i��$V= B�~���Hi��� l8��Yny&	w�e�΍'c�!�=�^&?B�"�mw�33�����i��s��g���%�2<�Wj�Z`u~���'�+D��-�q�4?��X��)�I���E-��i|�S%��+�r��`qs�P�vk} �J:�n��k�����[[�/��w�)�����9p�M�n��L�����2��WSl=	.~����&�(���>K[#�SO���]�q�<���L1	^rzg�"�țV|�Ӱ��#��'e�ʑ�?�K��u�a�ͤLҦ�8�7�����J���X�t��d0ʢT?�q�_$Ӊ��Kx�bRw��� ���&�N���G��tMW�<�5��U�;P��)F����b�*>&���il�cV2s���L;0��n�d%Qm�r������@�M��η,�4q��B�_~g�^\�	f��x�V���*�p�$���ʎ��Aq������/a�:�x׈gmEƔP���5�| Շs�̈Z$���zM	?�}y짧e�n���n�� ���HB��׹c^�]�*I�h5�.g[�Bwه��gu.��ivT����d<�0-�/�VuU ��C�?^����=?�'����'�[�����M�ͫ+������̒��{�nN�*A&��'������_�<s�l�}�K�M@A��o ���~�J��e�qB����^��=��y��M��ViB֝k�A���4��_���GS7�e円��<�>�>��{� !~1�H�`�_�(P�а9Υ�ٙ�9��t�J����n����B��è�o�TU��cu��Рgs���7]�QP�Q�訿�-���}g�����|�pSw�[W'�k-.�����I�瞦�.��G +�p�A�. �����}�oޛ �K�R�&���y<�����0kk��[/�D�*	-B@��0���>5�du���$�S~��/�*o��/5g�[�G��BhЭ�h�0�YJ?�tȲ����a�� ��U1qz0���D�$w�����<����.�]2Fy���_ZT�t�t�Au�Bg��oMS�q�������y��7���Zx��z�@��������νd�(�̼�pԢ�I�N�@��R���ɹّ���2�z�1w�2F�1z� �����	(M(���t�h=$�J�N�n�nad~�O����%h�����f7�B�ciQ�y}�adEr0��b��1]�؋�����D|�{[��$���*U6�rs��\#M�BA2C�c�o�\V:v�m�ў&IJJ�� zܔv`Z��j���;�y~��:H�S�ȍ8)=�n�5�q8&4�s��Y�?|w�+K�����ϝ*�V
���:�I�ѡa��F��'��%Z�"��,YY $Ȼ�'r�6�(�G��B���)�f�zv_Jό���w;�������F��%�ЗB�.-2���kNCQ��q
�_	'U���UA77O����8>TyOm�*���S֗��jA�P��-0��Z�F����QNH����\�ék��~��D��6��S��~ܳ�H�����0�p�,@��]$!y�O���R^��%�X3Et�X�l��XԞ��^9͞P*.��o����6o���<iR�4����o}�密2���1�B �-o��|үыjHb��A�T����c��]/�Y!��op�4��rE	k�I���\Ć�2S`���D5����$/��'����/�B�{M>����B����g�W$z�l
BD$8�1�:�Z�=��o���l�u�P��f��!9:�q���?_u���B-�mΛ��L|I�ܠo>��( �����4*���&TZ>�K��4�My�Īc��g�ʻ�xJ$~a������C������aBD�`כs��N���B��L2�y{VIT�,����t������eG�	JV#9
*�a�hG=�*��!�j�qs������-�!ۓ�wH�|wO�
5,Zd�6
&0~����ʅ�S
\��9_�?�&X������<w��uKM�6ۃ�=g��7j��ҝ�M$ 4V�4�F�D���[���Q�6t��'���\W�����;j����ѐ��wc�پP�׾O�8��MB#��J��f�j�j5dy�G��9˝f�س[��=��rݝ��HY�E�rt~��5�J���*1?G4_:*����������p���<��,�ou��Y��*\ �4!"vp�W��&��8#�V��(fm��l=%�~�PK��v����K��D�0{����ie�ת�<���eb����f �H��]��7e���g����GB��h����g�-Iƍ��[T�]�x�@[�R[�W����Sǻ�MoZ�&�7.�����N\�b�êUw�c=�rT��H��o��pKM�$!��ɲ�@��L/�ebv������-z�e� դ�!�J=�{qAq	X}4�Z��O���NDp�?���o�:bj~Ȑw�0��9[A<���fY��dY4�Ӕ#�zb��P�ypV�y�#a�̏��J��x��;����?k��I��R?/���ލ�POc��2T��=�&���9�)j<�1;�tj ��N�?���/�X�t?LR�y��7C_c������z�ʹp��L�ʌ�Ț������~�����C3ϺCe\ˁ`sn%u�xL�n�����Dx�fQ�};p��k��K�j������)1u��E[�����;��)��Zx����^�<�ѐ��E�kv+=S�q���d1�=a�ng�28�0�����	���8��>5���a�&�qL�.��7ޟpӵP(��3ӥ?+T<W�B��6)x9u��H�CK���°�u�6ܽ	��z�����+5�����>*[�ʾ��
���%��g1���y��s��%U�����<��Q�V��(�{~6wx��dόώ2��^[&s����C�Ky,��|p�����7?,Rˬ�g<m�gF��������n)�9h%�� q��_nU�66y���� �U�޻��е��93|��]>�A6O1͎�n�9e�Q��ez<އ��OE��3�kAXXT�o�2��9�~�OǸJ��W�{oy�N�KSML�!؉b=}��S���KE���џ��@�gȚR=n@�x�����]��{�{Κ��A,�>�&s��� ��O�7;�}��\����<��,��ȉ����D�j��9�x㣧��i����h\�����u"a��� �(��V��R�������1�.n�� @c�}?c���H����@ �������(�l>B��bPq��lg�툱+�8�����)K�R=�'9��K߅���wZ�B���T����J�>�xy71"��w11̂�7>�~$^_��j�BG4w��3��*RE�|ӈ�
���>�χH��b���^�Ւh��`��M�PQh���@�]ԗ��G�p5�p	�$y�D����sx75�P�(9!s�:P�|N%j;�@��|��,Dx�Ӏl��u~L�?�p�T�3Y���/V
��q����뾝X�Ϋ��exϸY�� �R'aQ�;;�Bl�&���g���6��,�۞�TSB���G�:wE=��i�����,�`ؐ�T,�#ۯ{�8���d����\>���ج�Up�b��>�ي��ؾ�)�38�w~V�GM,Q�=���S�.��um�Xvi_~�;`y�R����x@>�z---�!L����9��:@&W���r������O�i����t��Yg���E�AC���RNyN�.���Z�lY�][��aZE�!V��2$R2fJ���2�%��yC�
J����w]���sEP(	
Ձ�ɻb�J�a�q��zP���-Ň|��� ��;��Ѻ*�"�^���Fk���f� 
d��	�z9s�F(�\\\�"����PBv1(�=i���<�[['���h��X?!�`�a�<�nXn�?�+��gI�ob�ɲ�	Lg�Y6�����k��s�N7���6sc������+�v^n��!��"�������K�����F���	�����H.,$us�'���$��y-�$9��z/���t�u��e�K��,2�GZb�jn�_5���sRF�?X�ϟ����fR�;�*�L8�_Г>�w�\����ͩRx�pM��)��0h���]�<Y�B�N)0e>�� �sq�Cn&���b��9j�k�9���&,ӓŶu���#�?�Z�?)��P�+K�w�j�v����|�Y�Uk���:	��A4�]���2r(g� ���~�1;˩����)z�p�N̅�U4�=|��#�Ȍ�V��9)K.Ki�o�j��bS�����)��-���و��ʉk��lnŮ�[p.���)�T��ц:@���O��]@c��Y����������V�]*��-��8�)�Tio��K\�0���!�������}E��w��=�j"�W]�������?�<�y�(G�S})���9��6�&>Z\������&��J{=be\s����:Gs�X'{�F�^Nϥ���\�V�~=g<��w��}�����]��	F�Z�(Jם��"�c8)��w�Gq�.��۷fmEOWH\��5��<Dx��K���id�i�`v0ȐH~�����?��^k�fu?;�������5��;z�9��b��\����Ms�w��;N����Q���F���Z7�Nm1.�88m��E��ǭ�p� ��z\?N��csmqX��<���pԬG7�.
?��3�3�!/gý��F�)6<�B,����:�:�%���6��4;o~�q{۵|�����='�]e.�����[/B���F�����+�7�W����D��8z~��P�<"F�{r�E�L�^���?��,�"B[V��M���k{�Q|_v>�4�=Y
ן��K_2���G���⠹�����}�$�<�9NgrҜ>�|*[�8ⱗ���\����h��Y󉵰�BK{,�z
���\�����{X7�z�A��9G�-wU�)zF�֪����[���VG��n}�efu�Ё�;(��B��!r׹-���հ�\��s�+:!�,�*V��Z�N%����qxo
�hJ4�����z���L.���8]juGM��ŮL��Le�y;� O'J����~\�-�y҄�*kZ��XsXY�g���=��_dJ��i�E
�������<��6�r����r��T7xQPNFf�Ƕx��k�y|�~\>�{�%�}��9r���}t���V�413�;�Vvo/;��Ȉ|�	vV���Dma�	?�,�-pk��3)**�\�Wr�I�#U܋�{�Y0�GQ�K[[[?�>I�������j�Uk�m|�`��#ח�f ��q��]�ⶦ	��Z����t��_�IJ���#z����J�۶Y���� ���%w	0X[q��ȄSF��ԳW�"��x�'�
v���������{�w�4�x�t���Z+猴ܳF�}cw{r<�V�*3��`�h8����W��ӵh���sW�k�-��M=���Zv�+$�NR����j�rA�	Loc��
�Ə����(�;����D}���3k�Y�
kMp1�NY=llB^Sy�Ū4�en�E)���A��Ҩ�}�	q�kY���E��N]Lk�X�l$s�.<8::��(����=���K�C�������q��tT9M�"�*��1aĈ���G1/.|�cɩ&��kcm�[�X5�F���7p��+��\��t����7:oȟS�?T]n���'
(y����5�d4����ܖ��C�y���g�%��Gh� 6�2,k��۳����)��nذSF��K�x��,��H��\�� �.�l{�	��p���H�R�~n�����rlIRNG1h�7�sb�+��uH{���I��v� �de�`T���j�6n�����Ȥ��7_�܆4oA;Nw9���Wz܄��g�ٚK�Ӽ���y�Bu���e�$G�^4.�"��."b�%B��:������S�ݯIVs̽�iim�Ĝ��bBk�"[��O�1��o1�I�{�����aHwq��s|��-sG@�3�e����cL�����Q��05��u���N��.#P���3:{�����L<*����2zhХ߼N��!�F���\����x]����ɇ�|�A��Lm����cqB�V��bd�є�<$����$m�I���d?'����&���"j���`��1����OQ�K�`��\���%��M����s4���Ǥ���4Vc�ǵ--���r�+�Q�z��d���wA`�Ne@(�7ȑѡ���(۟%u������KZ'����Z~f��R��较B�x�s}�c�s�k�"wj7�J_Ǧ���.��/�kI��STId&|���9��u�J���f��\B�T���v�J�DAþ�yƤ��j� N&�ŝ�^j��NO��p�(w�{���tَ3^RCx!�������U��t� ���q�'�X �2p$���~��ӆhU�R��Ɛ*�O�efZ�t�W����i�4꨼=i��b��@k8�E"?���=<�*o$�N4��n{s��Q�mM���K����v�ræh����d3U��.�J�Y��A �aB�/�;�9t*�c��էMLW_���Z�@��n�95!*r��D]mm�|L:8�h��V�o�������-��~h���$�V�}���͌ڄ������ח!A%Y�1qH��"��rЫ��gl��S��Rp'���8FhI_ɍ����#���H����Y�׋���8�L0&��q��G�B���u�L�D���u(�������5~���7V*N{<���*I����8)J��4�r?ܶ�bL�IEY�W��woV�����]\Ȋf:E{8B���,8&D���݃�7�,��D����o�~����)u[.�)�c�M��4�K��"zB����:H�4YЋ4ϲ`N�����t����ͯݖ~*�z�<b��5�J��ɖ6��-��/RA��,��g��tw��d���o���S�L{e��������]��ZIp�<�&u�r[���Z��y�ڿϘ�
&�~��Q� ���.�۝2B�{�\��� ֖G��%u~��@�lrÞ���XI���×&qbP-��A��������V�(��[ac��p�+�"�ֱ$X�.�+>���)60�r�c����j�V�l{�Ԋ�$ ��<>�q�s#��:� �ͬ=�!����m�8���c�߬��_���?�t�#��j���~a����^��гB��;�i��v��?z�x#�ECM³syL���m%�C^��u��B�?���O>���Ů	W��0��n�E�wH��_f�t��
���.��>C�6���M^9dW�b�L�Ѭl��F���<N�܃�(�El�'bca?��a#	�"^5M�8ڥ�����8_�nv��E���!���7���l3����kK]�q���y Jje!��f�/���=����u�Y��"���#�F(ϲN��g�``�FX�"�A���|��孖��J�v���0�I��B��i���'}x�gX��E���h4ѡ�j�E���4o�O�rz��{�������@���r�3Q�)5Q m�ʊE�W�{3�V��[0Gq��0ԕ�a�R��̓
N����q';R�U�~g쫃C6f�GHG;��(�����Q�~W�.)�p����?_h�O~���E���`�3��ˎ���Q~1x��=~����$HLg#��zܞ��]�F�q������h����tꤨ"���^!2�7M�%1$�Y�Fʔ2š�����z��s��uB�}���6��qf�o�����:IDt��D�x��l��2_"���FV��*�����7�o��z�d�d_���j.�d���I$���"���?��J&�]����ڲ���uXGJ��j}��:&�ydV��6�QuM���Gx��BC�=l��(���-��hS��2���9�yD�̆�6I�͚�4���| ��P�ըOW�D�5��ߕ��OT	���Q�]�GW�悒�N�0�^hŽ���9����^�'!�������B�~oV[n���?g��*><��q~gE��ҥ�1{�WW�T�<�@+��ot�
�|��I2G[��Z���d�Li	G���c�:
'
3';���Z�$�>x�V�;�����| ����\h��lڞ�6D�9����R�����=ȎS77��e�jq2�Of��p��ޯ���;�d���o4}���K���G"�M�3.�{�a����=z�����F��}����8I������j�h�Ar䍻�����KS�Ompk���W��Ï��D6[�%ade���Q_���lZu1��E���]�l�����w��
��a1��؜C{k;�v���J}��Y��_ǡX�ѯw�$�����d�ū��B��g{��J|ۀ0���o�}QϜi3���Jo��a��!N��r�JD�DKR�|����V���Bq�D�Yֳ�jɚ'>����	iY��K�R0X����d��~|R�+��ڿO�%|��s���}ٚ=��y� �?��G�c�i������X�(M�p�e�f.{ؗ��(�ٰt��><_���]1,!0(����� �X��ٓA����?�Ur�=O������Wz5�nz�z.�@��v�5�]!�a	˗4��N�2��)JN��RO]TdO~�>\�A|�so�����4��Mq��,^��]8�>΢�f�����ǂ�$��s�E|�zm'�0�S�]4��g��7��@������l�K�ċt�'�v��ݶrd#��j.J��a�bv7���+��sr8��	u�����ڸ���1���y~@U����\6'ɏ�� ����Cw�s���0��5S�K�(yv�o�ML�}j)����e��+UAn�맫�ǜM�+[F��!;k������6*؟�`�p��B�L��*W��+�&��p�ϯ_�C�*����Tq��ClMt��-e�kϤS��1\T[fwgtu�c�GH�"�J�(:�C7���T��W${$�y���h���A(k�h�rB﮶f�A���矍Q�¨O%�a�1sa���`���c����?�um>��9\��;E��J��*�Ԅ�2� a٦��)R�'
k$v����e/��u��62r�"��P�:�Vs�	�FG$2QQ�Y�i�yr�BU$E:!��Q|f���:]|����s��f�����q���}�u|����,C������}zU�s	�\��9��m/J|*�����j��(6|���e�_�����Q��U�ϸ1O������_��Z�t�M����7��X"+�CR����s7�c,|�t�*�"�^���ǽ��X�K��l{�|8W���i�`��?6�rP6�u�c�6C-�?���7�.��υ!C��vm��	�B9sp�Z�b�q�'��� �����!�+�ytH;|l��*���һ�4)�N�w�ӱR'	����[���(ɛ�����z�K�O��?�@�`�t����'����>U�Sy]8{�ˍ�X@Y�]��ׇTmΰڊ�/�ܝE�y<s�Fv��c�=���)��- ^��9�b�e�� Y;��3�u�?u����|�(1s��<]t��Yg��_�i�O�]KV�,��"��7*d�5�?�o�Z�"C�{Mf�+�US��٧dh:��(ج����XA>����,�7���م�?TeN�I�G;_*!@\QKi,؇-7�l���w��ͦ��q�[H��u�P)��Y� �d�d�� �0�L�=�d�Ȟ��m�8�����r���~b���!!2���=������_�+!�g���oy�92~})����M��<�^F/�b.37������	������9�a����#Ł� m��Ϊ�(�E�8D\�S�U.��*����mۘ��т��N�$u�����ع3�y�P6@���)��om��ϫS�d���Hѕ�8�W��T����u��q�iw�U�QD�u-g������!�໷'&�����$t�g�~�r�l`S��w�f$�p
J3�F�g�녀�H�c�G������v^{���-n����rm`�������t��)s�쬎��xAL&��a�N���0>��̯������p���nVgK�t��%#D���Ƿ^_v����h�����/�J-�s���#�|r��X�{w����.��1��͟�h�W��z���e�d��M૸��]�uc�
�ɔ��Vp��u���֒���ЧJ�eɳ�h�������'���u;�0����Q�V���ΰ��	J�a[w������u��<ʱ�Sq�ʩ��(4"+����wg�DRl����U�`�;e���k�{���x�l�{�I���I'듨q;3_��7����鱒��4�(���j������!{=������%s`��KTug��-�{Rњ(�����p�=�����K�pX���j�qWA������&��Џ��Ct֫�~������h�<�s��9� �H�H.cnV��>.!� � {	7ec,Ó���al@�3'��R܉�;��������E,�b!"��X�ɛ���\-�o�j��Z������=<J���I] y����!YcG����9Ӳ_�ON�a [>V�X�L���+!��=�	�(U�:�p0�;CW�Ҫ��mz����V�n�(�7&����v���{Q����u�D�1�Cs���w��(O�C�c�^A�չ����?��;+7w�\�7oBE���\)�D��2%�s��n�5�A1�l��:
YZxA���c�Ղ<��7���ڊ�w��C�T�5����v^'�d�+l�]%O�sS��ս�P�ި90J����طB�N,�h�vɳ��K��L0�<�~u�>��y_@ό�5��$�����%���+4]�Ⱦ�݃R!��F���Ӿ�\�wD������6�����]�/�����17d�E� u������s����Ƀ���Ҽ�읍rJU�H"����1r+�ą(�8d���m������c$��͖+����D�¾��R�T�2����[�u݆+�LN�H�L��Jr�W�y�+���>&�gVZ}%?�>�z�\Dn`�N�2����!��A#��3���G����\�q�/��v�J�J�p������zȶ���u'�i�������Q��a�������j�z�u��}'�J]��l����[
YZr{m�+�]�h4r3U6ڱw2y�vny���	�Ő��X7֌p�<�����o�!{�r�tn��9X�`5���Qkv&)Y�����XA��: y?�A�o�,�,�3y7��1tE(�U\OM�E�[A�^
n,�����M�K�(>�P�Fz���Z�鋮y͏��5Lǘ�Z�8���T)7Y����O}%����F�60�_�3���V9��skS����g�m�D37f�-qmB��"ĆZ��_���.��"z����%랥Yi�.��^Ail�a����F}��իv���\;1v�e��L��o�!����Q��v��y��d筕�7�z?~y��&<|�{������Mw0��	$����M���Ȯj`_믁��FA�k�����3t�OA���e�(�w�;]y�Ӕ��c��{`692}���D]� J��,	 �DX˹3�f���9��N{f`�䌾>��-�������F�Ǒۻͧ)�{-±Q �����Z;+��rW����o�g�R��Nv���s� ��YK��A��w�*׫�����D?6��S�H��{��{�%d{+;��z9��m�t��U�jd��������-��K2'�����ٚ�p-]�nİ�����.C��㸯�6<�_=3�?O��Z���ע��ڕ*Œ�
=ht��r�-�m�w�p}�p��z-�p�CWeJ�j�B�����d`����ܓ��:qC]ݟ3[�����X�e4�o�oG^_ӓ�� ��s1-xݰӐ:pxprJ�� R�0�F��*%�q{�{�S�����uh}g�Zn��{g�O>6�hiߓ/��~�0\!�96c}i�������*�	�LW���t�?B�z��;q�Ĉ��~݀��\|4%�5���Y:�vԧ��s�Β�E���^��U�[ݐs,���>���v��@aY03@e��4U/�y��j��jb ��r&_�o�~v���|���*`�᪖�}��BV5�ǤK@�+��k�����58' � �9����d��pF8)�_�_'_�Zε��-�A����s�Ng��^b�O��Ԙ��^o__���lM�4\ː���M�D{��5��z��L�Z��^�����n]�O�{�}��`o�L$����5�`�W����E�H�G�?��z	e����|�(�h��	����(>cuG�HoQd?�A�����n�+���\C������������v��n���Y`�۟f���W�ep�'�RÒ�
j��>j�{b���f 
�U���N�Sb���Q<�T���@�k���F�QƧo�/�;��z�Q[P��j�&�>6ӽ	�A+��e]@O.N�h��` 
y����������p�� �ba6����%�ݔ��4��/E�ޚ�
�z��"���5���WjL2�˛ϊ��d5��\Dx��˂��a��1G�B{������T�H��j<��0�8D���4C��@�Ã�/���9�쥯��1����z�����q�%#�m���̜g\��:İʦVQӛ���w�*�%�	�Ś��ry yS�J��xD[J�^���Z����Kv��n���"�[=*�;��Sc�W����k9���~K��^�0k�O��ռ���1'��1�ҟ��Ő�J׬�l��k�ix�=:8�ŏ�_y|��&E�L,����(i]Ŝ�kߖ�䥩�ܶ�6s������;�� ���x�0��/������y��B�l����:�ɆQ=�Ō�f0w���,wm�"�r�)r�ss�KU%����!U�?�����_���zQR�L0�v�s{w�uڻ�%����������]D�jY��5m���Q�/�^�D�����(��>��S��ˠC��:V��]��e0m�,Y24R�#�㔉b��F�����h�G�yO
RD)����1�^��ॕ���k��.ׯm}���H����_�/"bQxm�JMIᗒ�nk�c���446q'L��1Ȓ��FΫ4�`��j1����+�S���Oa�L�M���P�Q���/���0�������R-U.!j���/E2����{�x�5%�`f3S܄��u��L���͛�<t��ggg�|���4V���]�t5T��!�k�A�νϝMv��u_)v��^���~>goP!܁JYu�(�)����[@=7�~�;f�s>��bv$��}��Ȕz�?�^�G|���#lT����X������1!b�U)D��ƛ݆�hE�0$�>�X�4Q\y�x�\���Y������ޜ0sC^(<(��˲~�n�FS��S��G+O�4;�{E�E���Y׃���"R�Y�ec����`��_�K�fu��Z�H�)R=�s�M������#����r��U�]3\sv�秳��z��إ
���-T�-���~��� 5L��[�o��/�����<�I�OGd���(�].xܺy?F��;��m�02�G��-�oaoA�Ӂ���w�ߍ�+#�n�����-"���]M��&|��!ZvhR�
[.^r'���N��Қ�����Qi� �^�������s��Wt}h9�Ӷ6�k�� <�#��3ٸh��������%�}5d LR�q���������r��o}*��W,\��:q�?�vK�$j�3v�9����"Q��_#�|a!��t��9��
�U{��_TT���,��~b�7���ˆ.;3����:h$�B�����tb>ӭv��vfS3��C2�P!�!���XqK��r:��7-Q[�/o9*�"w��ܝ3b'5R�����K�cm�5���9�_��:˄ֈӃu�3��u��~d&�rl|�`�b����Z��mKrwM�d��F,����mί�:�Z��-*�c������=O��ҟl��n5G&���k�O�i0ƕگo�R�����j]�fn��+�D�`��D��O�7��No�j�>�Mi���c��~���P�,{$�$G�Ǌ��lG�
��������Q�&78{�P�q��͝��{_���~���ǽ_���9^����K��k�r�R� 4F@�
�q�c6���e��j���`@�A��/�d Y�㈆�4x
�'_f�����+��ѷ��R���ܑԢr�Z-.���6ǻZ�w^j�+|�bjsg�I�� +"��٠1qgh~Y_$��w��=�lj>:#x�i�3����p�����
a=r����awF�!P�٢��Bi+��x�bd�z#`B�\t�X��U&?:m��djju�"�t�w��Uϭ� B������S�OvF���rNk+/oA,��o�7{�AU��v=F�)٘8>)��Wy�'"���W��eQ���6�堜&0��("����k�'�^=����m��^N�`�5��t.�ez�0}� �:�1�:��vM��q�`l?�z�3&���b
z27;�U�~�"t������wL7�	?c5��h�Ey�5���]�5�ps�q�[C�7�z-88�{@`��N��()��F,qᛰ_p�&�f��t����F?p�)۬�v^��%N�
.*���@=%���<��b[�C��w���(��[Q����ۃ{��8����5�nL}����ks��ppt[�U&�߇"BF�O:vUPg�	����m}
�=xx
��M߹���Y�0�{�]w�����'�@�xi%��^���3�>G��m[�\��6���������xT8cUd5"0)���OS�P��`OvΎ�����ي�56O��|x���9�Q��+bW��.�c�Z}����Ib���N۞��牄�y�U�RW�D���Ү�-�L��ɺ�67&	�
BwM��f�P�K#;�K#^T�.ff橄�׎yE���m붌���L�L�sH��;���Ҫ�G|�K��\���kB�M��j��/� �c%��͡���|�Z|�c�f�G�e)�<��p�������� ���[�%�r ��&��K|�tPI:�j9��}w�7���kH�{������ĕe���8AO��%}��x:�DRR�g��v��K�e��%4v-������(4>z\�#���r�bp���q���?�?2��cʭ;w�K�t���p>:F���ɪ)��4aq��G�D�/"JEg�F�5�`1O��u����2ɼh�\v���9_��
jw�,d\q�U�n��;� ˙)��CL��ΜivKл~����(�2x{,�<c�r�de�c����|��K?�M�f�S�l!����I�����х���_�U��N��~\)N0*e/#�}G���}���]�"Y�u��5�rR\�	l�u�ǡN�j?�5ߛę �`cs��U���xK���3�h���)/B&H��昂&A�NU�	��z�6��)��Y���X���JF��N�_*��Av%??���_1A�ߺkP�X�Y�]�*ZhR=����;�|S��EsƢ�8[���]�hp3�̯��f8S�Z'CW~��X`����fDF�����y��:?�#y�^�L�F�L�ɒ�~B���?�<����m�3Xkc�]6x�}v��' �:L�q�,�M7��^�*±�����)�mb�A��W
ȹ��0�(����Oޗ#��s�J������#Z�`z���A;�<6~�)F�*��ڜ�����$� �v���L/Ek�!e�Ҩ.{��ٷq_�B����	qa)|6�`ft�:iO�}�'%~>���� E����ű3�+���<����WY@��O�>��6.�Oz�7�H_��}��^��{�w[$����ڟ^�Vq�u��_�I�R�DF���kE��CQh|�����QL܃���(c>�B	s���+������ ^����܇Z��~�~4���S{`�E�(�#*t�Q��ʢ���^&�y���d#��El<
�i��xG�/�Z�0&b�_{�����U�1���h;�#&m{J-�Aޟ�,�M£�C��J.Z�1Ny
�8s��$5՞�@ϲ�]˅T������Ś�����(�V�ᜮOw������s`����|�n|~��7�`�8����cR���U����^j0_Z�TRZ��un����H�
���S��҆�k�)xa}H?OZ����f*��67 �ޙ.�B{y��x��r���:Ϗ>p`�!��:o�L��:����*QK�w�h�����[�_-q��U�!�HR�W� ��C�0޽�3���?�xN�4��.�����35�� 32�Ѝ��O�8�)�$NGV�\@�5����U������5�^�k����,��ٷ��~ʘ�5J[/��27&0��ǥ2��ON�+X��g=92B"¾s褂(�>^`�r��*Z���ǚ�|������$�ӨL�K%𶼾B���"�U�.�3�b4��tKw�Z�N�򭩈?������<�v�4���`���qm�Qz�\��z�����w�6kc����z;y���L�-���.��'KL�Ψ�8f��Y��Z�k��*6��������.����;��AmRW�3/58��O���q��$���V��&1q
$iM�W2�R0��V��1
���,>@��Z�s����g�/��E�·�*���=J(g?���#=b���)VJ����ˈ�z�nP��;��zqO�����U�������z����_(��1�٭�_�:O������?��t�3(�PB��.�?�@T�HD�&2c��R䂞R�*|~&�)��*h�\����߽�<�<"6T�����[}6M�E�`g����:`ܱg��9�ò�,�m7��ŔlP����u~7]$��L�<,����3!�BSZ���0r6�5�)�L7H�!:T��������gTA�P���CËY:�_
�Ҏ������x]�����,��)�/���WN~+~�+�$7�&�wvH$d)�̍�^�^��U�b]��&�p+����b��j]�v_S�,��=������"�K+����H�{<�l�ȳ��2�GS|ɫG�E��ڦ�k�nP���YlL����c%��޻TO�2����U �������J&�x�q���4;;c'���m�U?0�	�?A/m,���
'����
&æF�^��K���,���I��˅9|�#ٰm՗xȉ�=�J\�4�V�h���)�u�|�o��q�0��W��K���ޕ?Ыҷ�v�5�թj�u� c�b�6��^��_6��>�떨he�/Q��u��20:��.؟�[���o��qx�T���uP�#vǯt�Urs�B��X�n������<|��g��V���z���jp����/�� ��"� �͉_�Z�����H\���=U)#P����~Y��>��ű��n.m��i������c~aP�>T~�����"&D$C	hM�gS-	��%WG;��t�z����<K��*����y��������~4ӿ�W0���\B9��u�Wv�JDH���.n%�f)Bq�pw5�+��[�!��I�^�/�v$�o�ؒ��	�&ؤ�lT�C�8-��^�{`f�v��p�\��i4�d��z���\�d�����rt0�:/s�����!nY�G~���OJ��@ Y���{���L,>�b4+�������X�%b���>1�rD����%Te�ٽ������{
445模��/�C��L��R<��,*��)�%�u�%p�%�b�����:����A�I knOxnv+W�ݠ�<��;		r���v�ZdLV'i}n;�e���V����[$�F��Jˎ�l�q��e�LH`E����b���W,�x'L��[Ak�xy:����Z��n�⋾��Wz��f*�!�f)��t�c�����ܫ*9ε�]gˤf25ă�c��h/mK�{<�{��'��9�Z��:�9�:^{�솿0�$'MCIi���G��|&�8s���b>����l�޿�4�*#XJ��0���\uF#��=�[.�ӼW����ٜ�_y���c!0	��:��&��C�f����4�_:�����R�Q�!/0|&~��j�^ �K\z(��Ԓ���E)9E�?~3���*QK�P�E�.�3�/�2��`8��-�#9E�Kz~�g�� iIڮ�f��-��Wb
�uS�vj�
�XkO�X'ݻ����?�#��	 ���2=NN>c�Ab���~�_i,qbRe�e"J;V��d�J���e�.�o���ުI��7S�c�h443)��r++�u��&�p�ґf�5fJ-
w��KCo�AA2���0���t,y�z��t~Mn�\��ӽ���g�E��LGW@��e��۴�	CM�Z4�����&��~i��.��4�3֦�����86�X,�=9/zC	�^��<���2U�O���i�Ğ �����IX�^��]������l���M�E�~�h����G�ZP�T�׬����L(X*H��mQr5w��J�P���\H4�7����1N����L4�\���k�F�0����:�s�W��,��k�?�f��J7�П�Td���D�0�'��^A��2����w?���n�t1x%�VѶ`V���~�ʕ�{،�TTUZ�ku��g����E_�2�Ӹ{�C*�+I}����J#��ϑ����ɇD�*a�wp�>��q;=+�6��PSU� �{��L��M�a��'6�[y�T)�.�}�%N����)��(���A�4���[zf|���໘�A��7M�$��*��:8���y�*�%���uXu�WOȻ81�%'C#�Z�m��u�����~�]�p��
.J�S,⳵�U҅<Cb2Q��������bn٣��Ɵ��:6�9i�3e�S'�CDYbM��S9S�����1���I��وG�&[�V+�B�?�����A��pgB�v�>�Gƴ�Q�BnΚ0p����E�2��I������X �1m������adG��	��i�!��~�f\Ԭ��w����g}	?~z��]�8r^q5"��S������H���+�}�)�K�g�ӯG��M�W�Y�
�L�~p�}�j�;�U���(�7�\�C`�->˾��w���ƻ�`��o�E�i[t��D���P��Q[�7ӭ�$R�T-�g"PDm��$0�Ǐ}�R|z��W,�'ф��%=�$�rZ���6�B�d�G�ezQ��n�҇�>ɚ1נ���A����x����&�3�1�ͮ�y�%���n��u�Fw͔�rt�3[GRɄ��Y?�@����ٓ0�}\�d&��j�S6:0y��/�]��6����l�;�E<DוM��s,�O��(3���v��<O�����<`��<��mv�\���f�D���,�2�]>������<'��>�gee�x?���8�D[�
�9	;ji �c�<t�B����lUJƚ�R�/����jg���͈MT�!<;g���/@�A�Ģ���<CKɕ�gz8�T�f��IP�}Mbؿa�s���|I%4��Ϧw��Կ-/ȳpGݷ�������s��x�3Kk>�LZ�Ҽ�x�r�@��^���t]J��{v���P������L�P���xX}L�VQ�c'���`�}������3�a��O�����o��'�ՑRJ~í�@L��`�!�(5�B����d(װ��%�H�Zs�ʩS�i�(zL�̲F8�6�$��^�3������LNP{�6)�\�X��P�wF����ȁ���|��d�`��H��2��7��@H����|��8nHПB�|�k���A��� �nl����o�X+�q�*��-lvy)�GJ-�
�l,�r�6�[���S���ZS�z��^!7ЪlO_�ӈ)t��A��/ʞ����_��|$�;j_�F���Րj!��k،CH�H�c�+�r���i�T��P�嫻�c}���
�>iY���Q.t�7�u|��b���#-cp�kTϠn�,������Ծ���I
@�<h����}��go�D�a���kk�d��w6����q�����6�U�+o�FWG�a�]��ۛ��b��0��[2���>	�[�T� Ŀ��?�D�k�YzMV����v�9M�����Bt�𲊊�o�y.l��9g��V��Bg����n�K�%����ӣKŽ"�#>od�����X&o��[�Ք�T�&4��X�8#����/�F\�Hiw��_Hv�>]���������dm��;:B��.����A(eE�_�Z�2���P��xQ���v9W�]Ffk�
�1ͅ3T���(R�O�]#}��n���)�k�-�w��YC\"AK����<_��m��T���xBʥ�ndH���O~d��8qt�Q7����n���[��w�u���X���e�l��zJC�W��V�de��[�=n&$�����msF�O�[-�8]'�碔:�j杍b�g/f��"�4�t�kBc&|0�Z�#NS\���3ӶN�!*�/�9%�ۅ��յ������U��u����Q�e��	����,+r�h%�Z|�L
����e��Z��_ؠ�JT�Ko}wI��7W���		�W��X�Qq��~��Bnd"���s+5�~�0AK�SO���e�!�Bc�'�����Q�#�F"�n�lo�U:Ϙ������H���?�y��q����t!lS�9
q�\N2�?�_YW��$������Z8�����[����^�A�!��~(�f�ؤ$�Ms�2�b�p5�-M�O���-h�Sud��9�-�HX�����+�f�ip���;����;���'Hz2l��ى�K�nݜ�!�3:fO-Fc W�DbZ߷��!�W�m�.{
�ʮMQ.gr����߸������G�;>�(�H��KMO�/����:w�Zg�W�����d��,`����;�ԏ-޽�?p���`�Ǽ�wGGd�c=�?G�G[���������\s��>N��sM�
�U��7S2Q�~hL����w-Ż|�'�^(�n��͢>���VnU�r�H�_0����Z���s�z��Y���HF��'��f�*!Pj��戹Q���B�<������:=��A���Mۘ��������1��Q�p�(W�d�?0)�N}Y7��3ڻh_�,�]1�w/�S�O�1�y+:񼴊�9�ش��.@�m��\*e]����m���.i��@T�}o�DUF莖Y6���vp�H�����B�f�kQ6p4K��ZD,ېm���&,g�<��}�FG���I�O�����[���;����<#t�c\����S�t��hm�:ky��^0W���H�$�ΣΎ�����@�*�������I9J��8,�V���Y(#�_��#�P��~�Qw�Wֽ�-�:�cYgh��h��Hpl���\L^y��B����n��>Ș��$��'��7�8�j't�A���zA�x^$����g6�@����i�e�I�^���q��]��ǫ:c����UI+jQ���m�t���B8�����R������z&y�Z�0�Cjd�V{g�?=��.�q�TkSX���~I�":��]�����4���lUn�v�����~��B�g�̕��5�57�Z�fF7���VTk�3�,tqK��ܸc�}��xS��>��n�}>��H{3�����J���k��Oh��]}��D�d�ݎ�<=D^����D��,�I����<9�<وQ�>U�j�\6n�I��[4����`j�t�O7�ձr�|��j������P�M���ۻ��7���I,��ׯwI��|����2�܎ưX�Kم�o55/��&�� P_�~tTқ�jl�^f_�>�>���ע����S��4~�p�uM�{�+MKP��z��0�>6����^ŷ��{O�&���ϮlQ[�ڹ��ͺ��h���{���%X����^Z�ܨ��SEc�Y����q�Vj���ՌC��/,1e�dD�˙[+U+ˌ�A�����3X���_�ZҤX7��CZo�nD>ŭNp4=��/��UE�� +o��5vr�ן��3�O|irE�nmgNj�.n�z��@��x��S�C������X��)VcΣ��k�mn�jЀi�R�]�T��+&|��h�d��������\u�B<���;�vǬ�LS�K����OhR��~%�u�����'��)���L�����OLd�Ĝ|�_\WB%(��О���.�殛'On�1�>d/~U���:�}��y���	��z���(+֔M7Kǀ���/=W{v)|f���l�&��!���g�Q�q��ɵ��w�5��h���2�0�qb�h�V;��[v���^�w�v�KS��3���	���60��=�$�O���I�w��b<�}�,k��S�L� yUv����#��� ��a/�wV�M��2�`cG:X+�_�������PF����v-��p��Ȼ�N�$N`�n��Q8�;�A������=��\������}�MCC���F��_L▨��β���E� ���!����㎎�Bk$�5��`_�kaaa����@J��ɫ�������`aU?�Z��/���IR�l�k������P��p��{�n���[Ωa������u?�\��G�Jbe���M�z(��*�˖���5��LqeB<�,��/+��٧����	�������L���8$������o��Oq,I�vFu�LB��<�ݲ�@�_e�I��a�U͑���wզ�{��S#��;�캎���>k��o�F������w}�(�>���11μ�8{���
{�e]F��7�ag��X�"ʋ��s?
����_cyn}/����N ��g�Iq�����/����5�^Bl��ޛ׭�b>�ǟ�p�p���U���dMLpQ��JA�=���C�2���U��9�>�$�ײ�ob @g�R6�n�w��,���Խu��v�:�����=#(����7��|e���
�o=���:��I���1�G�#]4cS�y���̀:����+��ѶV��*�rn��i�%�^�[ �AEW��	V��:&^]N�1���l��Xκ�FO��>�V�~�ա77K�Q�,��7���րs���G�����*����1��v��U}s�H����	u��S������RiG��j���$X��LÙ�wD9�s$�?�T�xSj�޺�	K��~�7vav�����~b#��nŌ�u��������K�!���6�׺V#9�o��e��0c�>���']�u���\{l���������B}Y�k�AS��B��F3�ޖ�\)��Ҏ݋[��i��Y�5��=-�G���'Gʯ�9�s�eB�c�FK�K?x��I[N9Z�o7T�d[y���͵*��]9h<�K!���	�?�fF~E�Tp��s�ظ��X���;U\��Sv�7�7��ه���;z(p�KSn�����<�/W�m!w�y?��J�ȼ��v�����<��0�=��������dGњBCㅫ�%=&���:<}R��$N����l0RQv��眿ˏ�^i]��R��t��^�4�]��3	�K��u��)��ąg��y����Q���X	ON�'�w�"�g�:��FWVƐ[����Xb�yQ��ҩ���j�KV��D�ڌ�΅ɭɆڙ�W��6�pZK.��ry�p[�[��*�eLT�n��np��*������µ^���?N��岒�!���%[
�����\�{yC�?��R����L���]��O�U%�Y����g6�.")�aU���m�^��K��F$�����p���������Mc"<O�ɸ��:{�9�*{��w�b�x��<�)╩�����!���(Og�<���aE��]�0JS����%oF�`��o8(Z|u��#ా��6�R�8�LMM��Y���[�mlX����['UoE�5\��=2�e3e���:1v��c�3:�����ks1IC̠�*�8�ޘP2�g�kФ���M�Ԑ��v�t�tRu8��Nlm�n������F����΢��N4#���B͵��~�!:�����f:h�2Qw��|�'������i9;�h[CI�����q��ӈl��}����M�z���H��*��u����H��brn���;�~�����+�̋(���<��4��Dy�qǎd�
��-�u�z;���'_����i%@I��p����T.E�Y_����#/|�G��+ꎫ�.zډ�N��-�-��'�#N�ǆ����}IWt᣸���*������[3ʃfd���«��iae��
t 9�|�	<���ã[��,<���.�.�5����7;�N�]"����<�N�?��V%:^�U��1a܇>�k�� cBr��3jnH����E(��]<�[�°.�J�o�Nxa�r�V�ت򆠡��߰��u��
x��[=�D�'��GGzt� ��>{���<���O8�-Ğٷ��Ϊ�yK�h�Cj��X��7;/n���(��x;L���  ).�kŬ��%[V7��͢q�@�Ѯ�R.�A���kllM��$>N֗�a�G�'��'�����������Rc�Q��)�; \[�l������zK�4�%>t�l]}U���l����5��b�=���H�t�E qg�Ýu��hc��6>ԏ>JD��o�X����8ʨ4�����[�*�D��\����\�B|ڿ+���)Gue���_��Ǘ��9���(g��d��#QW0E�@�{p���m����.e_�?�Ԯ�<̾׎	>*�c��aqy}��$vi���1
��0���V�ޝ�C��ЙO��s��]���LqIm�dۆ�UD�Tu�po�_��dF݄CY���%��{����������ki����Ķܛ�8���m��{V�3b�u�r�N�������zM��dz��$�͠��%JZ򺤅S�� \�m46lK�]���A���&�%��_\���e#�D�n���F���m�~��P�M�)�b1��������&J_���Dr�->oo1�<#.b�q� ���f�E��b�0e�8�\����;�Q*��%O�v�����aS�"o0D� j$s�/�}}B�����Y�	���_�ћ�Ï������}�D�PȐ�i�m�T}����&%4O�!B@�/�{�%�3�D�����
!��� ��0�xf�����	���J8�<�|����NA�+�ؚ��g����Ͻ�����:6�׀�mu�m�j�#�T���;_9�x�����P�-�jh�!����뒻�X�A����I#CY���]�%�B��1UJ4\Z�c���Ո8��"�$��sgy�_h�4��U�&��ϊ��|�P+�����͇\�F<�ے�?��EN�sQJu�t"d��d`�qsrОk������.}�.&�;�&�(*v;_����n�Ϡ��%!7���*3���F$�	ߏ]���29��?��B7��՟}۵�W>���������:�)��eYdy�'�G��Z�Q·������w���ƴZ])
�oݵ�Q�z�6t��oߘbۑ������O�ֿ$��l�-8�{_eo���vx|�(kM	��'�]�\0�ǍjL$%���]��T�cQ6NF����\+�w�-g�x�_r��`�fG��l��߆n�'dU&�a��ٽZciI�J���Jۂ�Ș>�]�C���t)^��sjs/��"M$�5�(Ux/ɱq\S+XELMP�n�|9m.�\����-�f�+ rw)7�z�;[Dd$tu�T�6�/��Wڇ�(��i0(X��|����/b�a�g�Ӥ�^����U�G���L:z��ç^�>���3k0����
�� ���%��F����!
M�?FЏ���+�/ɫE�ql�<��4�o� :�2n�W��H$\xX>T{���˼ǿ{`�>40����\�fD����HL��<��=�sz(���MK!�s���vaycK�f�.�据�S��
�{����hm��Hܺt��]Ϥɿa��@�(���Ӆf�Z���ǭ2n
j~�;#q�$���D�}<�{g]�"j�r?K�`�x�~8���"�\����
��bL������w�������x�L^l`����nc7��|/����>�\�܌�K/t�W���W2�x����ݬ2%P����1��&�P��˷-�cy���ê��&a��"�lO�Ѯr�m�Ye�-�HTR;̝����0�k��eC�|��҈�q��<��P��p�������a)����=�����\��5gW;��I�x��oPo{�|�U:?��I��=0��}�ECp�b��u�bɀ3�&Y���;��z�������xN���O����OpD<���P�|�9�I3+��4b���j�[��%�8#R��%�  C�,Qn*~�AvMM�RRU���^^2�u�9񎆄�	q��/j�#��EQ�o��:��SA~[��1�Tt\Z8�i�J�Ã�+jjs��Y{��c�W0�r�Z����oN�e�������h��k���/>>K��f!5*��k�`�PI������Ơ���u��C7=]o�O�C�l �B���^���lr�I%N��W,.k��kPRg�
����^O��㝈�3>X���q^�B�Ux�͘����U�>
�����h�k�z�k�Œ���S{q/�,�����a������:�1�AH�b�S���-��W�erNghNWn~ј����;�X�.;�r֐,gIr���O�Z+#`��!Vn�8م�fg2���������%e%���|oƋ;/��R&�X,�=E���r������$��<���s��{�'h�2g}<�����6 $��Oj>���:�������׆[��1�~�� �$��,ʪ���[���<���ݚR��:9�����m�'��r�8Y�HJ�ƾ�\n�q\�8�#k�Qh�֍D�.�BN�rX=E�$~��-]{�L:à8J���Nk�Ew�ID�%�0v��g��;�����J�lw!�M��#��� :�s���E�;�g�mW�5��뭜�|��kG��+s)H�+���<��:����*��p׋ڤ���h���%9�:?6A�Y�|!v��}��v��^=�����7��:@9h�Z#_��<%��Qg%��(�ԭ�*j�sP��o���o.��'8��'̷ߘ��0��e������-����V5���> *166��ge}�#,,�́���<y�9��z>�IȚ�m�9F  �J>_�M�TC�3�+��a�;[H�s@���7��e��T�r�P����/�����rU"�h^� ƭB�ؽ��簀����S�ɝ>w6�0���:�K*\o�e���>����2�	%�G0��ҍ�?t���Q&�N}����1L��Ŧ����T���ᆚ�L>����^?���2��_j��i�߫N>���/�N�x�uv�V�NA�g+��{]��� ����u7��3���t���I��&L���.��������`��/m-�a�%=�큡�8o�뵻�a���㑬�@י��&iiIh�^X���OVso44�%��M��2F^ |zrlp��"=���pJ
v[��N�t�0j��M��f�0����� �W�Ltv[�!���).�ɚ�n�	۴*��[�+"��v�1SI�L��ص�ʯ��&8-�S$���7_�6�t��Ӏ���Wy5^��\�2���*v7�/���?�h8��������byw���I�΂��v�	ֶ|̈́j���MYgb{u����U�~!%)��Y��t�y���� ��5�Ny�'݃qq���z�5P�4�4=�5	 SBئ��/��aEWF�_��i߂2tm���:7�sff�]�,|�����-cšt	X8~�����Cw?���QF8U����L��J��$����O:�-��e��4疤��У(�J���1�df��	�v0N}�,�VWp�|�ݢoi�@�iQ�8]F$��S�b���<����]�����dU)����1|�1ǤJdd�I��aУ�����M"��C��L�V��{�e�D����ƶ�Ł?�D�u# �#�w���Hۦ�û/��$��Ia�h��6}qN���+i���A���� ;=mqQC��+��~�Q.�S:��W���­n���%�1םlp�����C������q���" �齖81���/�(��Ay� �}��w�G�!QQK3��f�bͩo#��;��n�W�5na�<��l�>�{aռ^��8܌�'nXO����cN�/��w� י�h�)hc����$��Q�i�G.�1G�j����KS�]ryE���ۋ��m{h������+Jd���h���C�i}�G�ZR\��+�ܙ�+���r�9���r#0YC!&]��W˰?�K�]L8V#h4Cjˎ78��N���3�7�F��7�&M`�D�3x�&K5����O\�B|ef�|��qS{�5ccIeݙ;o�gbV�o��bŜ�3�!տ٩u�	��P'��y�ߪ���XO��;����
�<���Ӱ@��l��}����ON蠒Y9!"����4���r}���B��{%�<�Dֹ	q�����5�l����m��i�?}b�=u���ϡ16f[�艔7���1ۙ�ƙ�޺3�n�71}c��ڙp��* d3�{A�]N�w$�t��!~���=H�t@ۨx�����`Wr���{��z��8��8]����?����ȷ1s�
��V�VFk�[0<T�0I��*g�z+r2 ��I����%��4#�8N��\R�����K�Z��/D!�;f�$M�\P!!a�ЄT>�Ȃ���{Zg������z�m��ڌOO��-ʓ��*Ch�����=�[��Z�HN�'0�d1?k���F��;ߍ�ݕ�bv��SPF:�af���oYZ!@ȊJ�Y%Fά�v� ͤ�n����x���_< �kĵ�\���/�9V�Ky��o�z�����wOS������o��3�Vi�������'��������G c֬�+�sqW�к�D5��n�e݇��o9�7���\9:�������$���<�Nh��o���C�^���� o�x�݌r�Y���ַ�g��K;���s�,&i��i��L�D��=3�w�F;�ϔ]O[���>�!<f\/��'ػ���o͑tA�-��h�6��x�/[>�wvA}���ge�p'K$T)�C�,>oJY�K#a8g���h���e:o����]�����Ŕ��JT���8����H: �ڞV~ϛ�;p���n x���&G�����������"1}���Nv��Q�����kyt�4S��<c']���5nn�;�W/[df�����3��R��^���+��� �0�	(��E,qR��ٝ�pz�Ү�
pX;l��&�(s SG��� &�=�;��P�9�7�+�8���ªV_�VP0�2}ǙR��8����H����[E\*�l�l���_n�פ�A7%���㫞����g_}�]��1~�����	�� ��}�Xb!�&����NDo�����7��X����;�~��A����"^�mk��e�?�X�碌����98�By�?�b�g��1��s��v�6��a��-^rh ��>!�RF�"@�Tj\���. 6.ކ��S��a���i�@��DV���~��g/��n$��<P��y�q����}p�J�K��u�AE���VX(��"΂~1��1�yf�>HDAx���l�$Df�,*�%*Jk"��e2G���3�	5���1�����*��e�x�=�׻hD�74�ԇ�<�C��2�B�ԋ�@�]�M볁�4�In;q���t[w2 4@�(eF���>=@9^�,_�{��M߃�O���y�Ω2�C��W�s���5��~��
ķ>]�I!��	��a��D��V�t�R]%�Wh�`�'�AkD�l�#c⹻e�\NS��2�+Q�M�
wL�lB�γJX��Һ�[�)�@��R�Z�>�L]�U\F�fF(_��D�m��5�s�:u�qq�)l�5�9AR��#o�A�����tϸ������0�Ah���<̡��T�$B����/�%�煡��������'[ܰL	����	\Jy	��n+Q\�?��g]ol��[�Y)J�\�hF��d���	�g�mD'�G�{xٝ���vN��_J2�����\|0ש��ԓ�w�`ΐ��㞧�%�1�|�jm����@�_Ƹ �[��C$E{�=�57^//�R|6r�a2�ϋ+-
� ��F��	-���i����P�b;/��W��6��㹔#���:Ƀp9 ͒����0Fmf�ώ"􆈐1�̡�[n���e�5Q%��
��9�=x�e�.���IA��Ǳ܆uwK膣Ezd��a�w�l�={��YӍ��>L2�z�xl�|D��i����%,��kv�QG��t���n��J)����`��l�n8e�Ϻk�'|��ځG��|G^[Ա���L���އ��x���m4��(r�xU$��O��A���8'�ثD����k��?@҂Y_h<�!4�Ɨ]�/V�+g���>�4J���J�}�x�VPF8c���±zA��̋M��g�|d��d����~FiL��cA�j��%�@>c:�+��Fk�0{�,.�ֶi^� �(y����>p�sSx�=;;���yѿ3[+X�qo�Hql^�[o�gvGN�uM�/��f}���Is��F�*-S˟F�}�H�k{�}a��`"�d��OT����3��A�hy	O�;g��ZlS@�D��Q���;%bo�6ƞ��hg#E�U_��F�A�tH7�)
H)�).H��(]��t�t#���� -Ͳ�t.������;�2���>���|��y^N�:>�?�+�mi�|��eA>TߠT��~0??�̟�o�~�	��~�>�������d�;]���W=���w����Vɳ�zKs�_�F�,~"`S��u�kRA����4�5>���%	��_���~b9�+0_u4�:8�h!w\������c�졏��'�e]L?K\��5���vN[<�u��H���ʍ���{�gU�L���b�PD�#V�	�9j1�F�|���qv̛���u˪��Of��fQ-Q3�)����QJ�T�5�t�lR�]D�`qÝ_�Vۗ�O���,n��X4���u���	h���O&	:e����JZ�$al�}g�H�#iQ��@��3I�����F���&�7�lFq�	g�5j�Ky��1�&�z"����
Oz��^(x8�%� ����+�M���%lm�}��N��w�ҍtw����r�C�/�q��̖��Gs���`G�k�u�!)�V�z4�����j�%��+�д��f��/���j��K��w�����nj�l���ߴ�����+�W�x���2/�p�r|�=a�b��'��g�����*������d����o*�d���x����f�ec�
`0F@���]�_cZ�i����=<���$�	��>l+}����7}�u�퓍�U��(�.�OO؞����0ER/�`�0^G��,���Oz=!o�X1��r�z�g	��ڊ\�����*k��K/K���/�g8�����{�./O��O��`n�&M�ۃ�+W��ʬI����B�0� n��+�
ד�F���ʌ	*�~��3O�/�G�J	�1X�-�����A��nͼc�zXF�i�7�C2�/e�6���N���#�6ǸfS&�_9K2*���9��PU� ����pA	��oO��
�6wB7��xK���3�TjĊ#��0y�H#*�[����.�V��v]�x�>r�Ű�w,L%���G������*wh�QĜ��i`vl�ߛg�k$�=	o{�֝��eo&=�.�g&�Ұ�l�lﷵ(/���4��+O�0l�Rݥ��`��$S�V�<�LtҁtWJ!�f�9�o�������bf�u�&��kjK뉢�̡L/Z���0;��L��������+שmwZ�2���4xl�;)�8{e�'j ��ۣ�M���:=�.T�Ѐ��H��0�.��������1ܗ�L��ó�?�/�F;׍��J�iᗕ͠�M�
��-��J��	 � ��1J����ܢ��NJ%Ծ��4M��`!�>�>⨞u~қ�)��S���V@tt����:��'%%7촋F׷�F���}Q~@W��٠�lXǏ�A�Ȝ��j.�Q�'��y�����'%%a`t)���	RNz�1���?n�>��*v��b>��� �/��1������K���l���p}���r�MҪ��؛�-{�9�R��S��﬎��Xzׯ_�5]rH$r\��֜Q���v"--��2�Z���}P+n�&�=�U�bV�}ʫ��yN�7��zh3�O
�Z.�:��̗�Gmٔ=�D��o\c����3�4���18��;����o��?�`��>�>���B�s�(�]����ǃHܦN]$��R���	�!Ѓ�RD�G�/q5k��z�$�L��zj�3�5�t�%**ՠ�}�ֱ��8"˞�c�Joo���`8]r�E�� �v�e,t3B�sn���\Џfu��ҨX��9�0��>=q�Oc��7��/�(��j?r�������I`� 3L
��Sϱzܵ�>n�
 ���'ω~h�9K����$��yм���U�e^s	����,�b��u�+�G�Rn�<A�m+�F�V�3R2�9D�:��̇�������桁�\�G=#��R^jglKn���w`խ���+����w�^[y|�(�SU����������6�����+���er����7�.�&�m4�wu�5M�^� v�I�((��}�ޣ\���=n�)���-�L#�h�dۋG?\����4�4O������
�	�*s|Q����9��J��~:��^��ߟ�Z���$G�G��]��Z�.3�E�_`����O���,�PN$=��,��4P��y��u�K�~�;(�|m2��|!qT�!_	�gy{7�� �^:�1{`�J7!:��'��\T�zA��İ�����/�N��*�j!�&��xG栗RP��=�=#�aΣ�W	J�۫NT���Y�z���hr'/It�J���T�{����u��@j|�;��N��b��S��?�ң�?8��f0g��t���%�d�s�$*����ћU���B���٭��?����5���uӼ��ʀ��r���W�Ύ#9&��ݗ��]�ß(Te���^���qG�E`T�Ys�Ik�Pgp���B�L�rt`z�g�h༖������ך����3Skf�ד+�g�M:rHZ���l��'sxyw�5��< �d�&br��/���x�߈S��Ⱥ��Q�g����JK��CV�V��)��e�u*�҅�02�a�[0����c�n��hz�|(��@�9�/��^X0=��%���x������.a����m��UQ��&0��?�[�yy��� ����	fMϵ�ټ��<ݩ����]8�Z����������fD#���I؁�ɺ���8+nӆ7�X����α z����D��yL����L���ͪ��S���� ��������(2NAQ��#_,���Z1=e%��;�QPS�ۯo�@֤^���Sֆ�&l�(�+�O����hf�W1t�J�������SW��-�]����_4Н�a������"��/�;;Y�C��4��0CTf�-���-%��L����ϊ�`�.���I���G򀿖N�>V��gK&����4mx�x�j���.��5p�J�^�)帯�A�1Pm�?�	��QjP�֫���ο1�4x���|�?�d��&�V��cA�M�IR������)����f��ͫWM.	/)�<znӭH�uuuj��[x�����OA�WC���˽_ ���lf�bIX<�_~��
��������t�)�b�T7��ñG>�{~s7}�1��b����W(�+˿["8Iq��h���	j����n�����@M�/��c��9�*"}�/��jS~P�8�{���r��o��
�K��^���ٞv�K�Z�׎���(�����	$�ڟ��6�_$������	8��TZ�d��z,6Y蘿��	�#������kX�BЗ@��g����=_�0˩�p�KJB"y�/����D| �f���u�sj���t��s)�7��U(:�֪֡f��ww���M��l��?���U�>��R=�~x�zG��W��~�d�e�ե���s���6���y��p���d\=QB�_B�d#�L��3��]2m&�i;~��2Iqѭ˴�D$$p�����i�&UC3���.6��Z�!�હ���+�v~�X��o���O�N �P��K����$��&S�ne��25/�v�$�q��az��ʾ�d8eU /�iT<��bmt�%H�M�����Ә�p%oP���k�|�8���m����qS�4H��^��bLb�2��Tط�nX����?�u���z\�Pe��U�<�Ү}��DZ���C?v�*!��4̢t~j���E��O�?���2tG�F?f�T�avW&��\%��B6q_W�L_���B�ޢ���ۈo�vj��X���2
�u�x��g��ҵ�ǷL�C�sS������q����8��|	.�mX���}�D�u��Y���mʃ�K��[2�d��>���;z�J�����?7;�%�htf��y�j%����=Ce����E�0ڳ�clek|��J��b#�m��ҹ�����A��]��C�[��sD7��j��;�)H��^oMb�����Z��w�U�x��Ȅ�fP@`1;�L}��mp7�A�����:Qx�9~��i�8tvLH�˔���t�P�� ��)���Y�㍝�S��ț�N"Moӛw���ulm�"��>k�x��AgOlpr����I�;��u}�w!\*c���.�(~SV)1�����������t�O�V�a���`��8�����,9�+����z����sA"}K�n<pd}?���Rz��!�&�t���b������So�ĢP~���ë>$c��M[�R����=���k��'���G�`�bg�����\i����B���Dڂyn�R��2K�Ϗ��Vwn�����2b�a+�`uˮ�o�$H��������ӾR�ܱ�D���$��%��G<�R�fj-���X�-�RJm�H��{��8��XI�$qj)9�A�/�~+�(y\2Be��=��@�5O��J���/�9$wq`�{�-����^���0�vzv6�{{��+�I�[�rE	�y�s�Z�G7�z�$�[CXgwQ)��C�b���B�����P�u�%Fq�Ge����)��usV|�eCRB-n
Ov�ަ#���y'O�}��	]v����%a;CD>�S��[��3�RN�!	$�:����XR5�\vI\�t�/��*��A]��<��}��Ŭݞe@���_Cg��l����]m���Z��YA2�9:hZ�$g��R�47��5��(.�@�XtJ
~��m.���s龺ݹ��$5���\J�1�Ҽ#`����n�K�V�Mq"�X<�V�9�8��n��/D��6r?��J��gV8޶�V�T�z������"[lf,�'G�����U�����Խ%jo0k��@��hM�"��Na3��s�o�x����a���1�&�vv.05;{�	o��q�r���Xս�7aByF�\�W/�Z��vv�|�C�(K��ڸGts����Z����0�c����as�}]0g����	�{�@��KM��l���lr�1rx����6��e�r�JL.Ԯ!�PBϩUpxTi�?����_�*B1��_"^���~�2��fO� ��h�~�.�����8�쵺=���V�K�6Oe�%�e���(I�#���t�t�!)��"@W��oN�6��Do�/��J��o�B�,��W��gBKʘ2�Y��<O���/�̓�����Ѭ��� �_[�k|ef��;�o� E��]o��2r���^����y�߁z����kh�~W�}�LwG�݋ɞ�M����^D�9�M����k�_����~Ҏ#+w6�(1ѿ�]����+��d���Q��L�X<��Um�/
w[4(��CR�t�@L���f�.|o��VO�A�6K�IG%\���Df������ck��)_*����4�{���k?���j��NrЏC�%�o:��(�xH}��fX�:��I]�Z���sN޾�:�����������o�LDtW���r���;e控\�wk��X���l���w��l�����$-����v�;�J�BW��!4���H�S5��s~/���vg-(�^eċF@I�6�NfȞ�l�>�>�kd��9����z)�������JEOO�{C�y��ig�6¼���rglt�I�ުZ��n]E:\�3�<�j���6�s��W���I��M�qK�"����e90����W����c\LD��g}���H��=�`O���o����)f���96v�S�ۅ��%�>$��-~�?-5��1��E�$��ޡ�&�8��9���ou2<��U�lݔiH�����cz�=	�K���c���'��d'E�F+�WM7�0*iկt�I�[T3C*��~�	p1���s��v'�_�|�u�:�Y���u�B��T��T�k}���Q�O��:s�����
r��w��)�wf"�^E!�C|�&��B�J� .��.�}\X���tB1�៙��f��W�L��U���*wPki=*�3���q�i��)�rN`m"��3�$^3��X�d�����o��n���<�����x��,h>t���� MT`�W���0%gp|���Ԓ!F��}�ao� Z�^!�Zx�p��-�fM�U�E#(�����˦`����&)��沌�K4�h�,{~d�ϫGߍ������K�m�^NVA3>����D-����Sծ����'y���������([��88h3�h��`@lH�o�k�P�шG�@U�y���k2���U�D �lȓл3��,�!���������ZR�E�-z1�_NT��؎��De���,5�$�����z:�g�z8����į����G��j�'�tuu#�8B��p4G�f1m��ނb5oW���s:Sc�Fm�|�D��эT��^N�Laʣ��H�x��є7�u>eh`�j4� !T񋋨ܢ��%�������C_���)���jC�+�J��z��bk���H$>�wû�➸,Z�x���K.�lV��D�� j���W�BE�6~�e���Ncͧ���Ks8xj"�KՈ�w52�
x�&6���yl�P���ow^�I%X�#�h��ݨ��W�B?�͘m���pOPH��+6�����L�7��[n�Td��)��C�௦���3:���/}�Ĥ�^��!���,7�譀�E�e�#g�̯I���.���S��6���5�c�<K$��0mI9#u�����?C�ȶ�٣�B� �m�����\���Ob�wIȊ���L��+(�dw߱���1���ߝ������0�r�n/{N`��s��r�~afV!E|%0P�L���+�o+$���I}4�mv��9\�J5~jB�vk��q��;�?X���ᩒ9/�ð~H�7�((�6�6w�����W�'�s��	���Iț�?�7�B�T��8���o	}7yҏ�_�qR3 ފ��poC����sΤ1��E�x���8%d��T�Q�[B߈��tW��8e���	]����iS�I�� �Sv��U�Y�$��5��0?T�
I����^��UA��^B���K��׸��R��c��K46��Kw��4��`�+�
��'����튍�8���t��N�4Se{�0���&�^����8�ק\��EBe��0�����,��!����
Ǝ��\B!���&�!�X�4�zw���>�|��3ڬJ��H�-s���g�/���=��}Z1������|Qbb�]�k����ڡ��|���N#��+wr?�
�i�����`��$x@��!�mEg���1�,Q��f�1�dswY��.�an�'\�;b�,Sh�dG5FPL��v���0 ��H	WVV�Z���[5�p�L,L���Q\�'=YIH�����wk�kD�n�<����L�j���C�.ںl���ġ�UvP�Xp�s ˩���qB?��� Ōf���`����6��^S�oꪒ������h�P�\�鿼���;���f��
�s�����}���y�PyѪ�.y�������N�i�+�Mxk��w�<߯j3C<]<��O�p� ���A=��<��ތ12�(���W!����h<d��Ӽ��.�̭�g�?�Hgc҂�ؙ����d垝��K�sʬ����)�rf6!M?/��3|�g�w<쩤�"1Y�̨�!�������@P�ʱ�$��}das�2���Wפ�w�M?E˿ҿ�a:�4�ů�/��L,�����G+�-7�@/�~2�ؒS>�Ǧ������;c�=��Lݓ�. ��"�ܦh�J�A�d}-͔�ʔ�k�yF_�l��DRٺ�G�3������1#vc�� �8��^�6=��8m�.A
�4oY9-����q�_���l~��:���k�� �1�_i�|�/.���"��Ռ�?�c�}���p������_O�x����!�6K��5wqQ�5��<���/)���2$%L+��������ء���L���RM�޸��g)����?>zA����������r��m��KL�c�&<��s)`݆���.��r���6mI	5i�D��4�_���o��x	�bO��ʯ�av��T �	?`�c�?�$K����KD�ۇ�a=���yRm9�7�i,���n��oO7�j��Y-gH�o)K��D&�q����#P�f�?��L���Q����C���}�7��$\��ր�ш���S���,���J��oʸ$�g3�ŏeԌ���}��Ny�����/h�HiU]ޥ�W�Na���`պ��o�3�2���]l�/�6"���V��D����o��z�����Ï'��<�)4l�
n��{H���Ҳ�+nm�^I�?����<>R���}N �
xǧ]e{'в�U�z��ן)M���+kt*�
#�5����� I# *��:�L�m��#��(����)jH��z܆R12�D�-��y Udx�cI�� ���6ZA7�s��\����/�!�p�=Mf+�9h0[2��-��u8�y �AbT>G����Fx!(㾡ߠ�`#`��[�)1�p���̦���-o�ct§`O��YT`��GTM��C棞|�򋷵�0pQ*`t&�65�T�w��I����9��B�����I
=U�;6x3O)�v�����cD&���כ�ұ���5���r�z��l7��s/3�r�J��0�<������������"TC�"'�p6�f����(z�q��m�N�;�-���/�a��W�����I��t�pf�HQh'��*�2��%���"f���;���������q��J�	`,WJG#����RO"s4���"�/H��Yl���8�������("�KbY�{�ۛi����a�����]�|ӆ���ndd��~'�!��D�ˌU[��ޔ�8���8��Z64d]���fH��S�D�����J1P$�`u��5��H ��F" RS9���IQ��.�Q�砬�2�:B��-�ȃ�s���ܾ�K���T��x���+Aw6᲍ݭΘ�!@Ʒ����"Z�}�rM�@�]Z��Y2h���٩A���O<���!�S�d�Ƕ4y��##8g���<j~�f7S������C���5X�Ϟ�Ȳ�ʝ�g ��&w�����N�5�X���lܯv��X0��M��-9�}yԫ���&ɦ���T&Џ���x�î6�	��hۼz��\��T�#"�xҭK���M�gI��p�Ͽ��9��Q++��B!�"��M���|�b��h�*O�J��f��ު}}u��Y�@�M�!##P��]�b@�um���O���DT�FKG��*�VH��|�L�=�نm),:�5l�E.�L�7!��v�������vM�ߩ�c�S@ޜ���-,:�MQ"B$���@�jo����DG� C}��Ϟ=s��.Y�t�ś��ݑ���e��;�O�x~���K��y�x��~"�30�k�e�[�$���(�_�--M*�pH�����e烏7 6�����,v9G\�{H
tJJ�D`�"�W�ؙ����Եy$�;�&=���B���A1���CNa[��"�s��u��}l��2�,�C߻<ȁ�����|�s�>���B�_Bߛ��W�BNr{��Kn��v�zV��`�@�$Ӟ|���90�j�&��F9x�[�D
'I�S��|RS~��N�;p�>kǳ���fj�����lѧy��vl���
��q�G��|m����ǂ��̬%�t0o���۸P�<������p���MyQ�p�^��V��M����pKy��'M1��A��������صq�٘���Om�ޚ���?��b%K��ӆ�U+�d��O���Y������Ŧb3D��L�����FT�3W)���̮o<��c�
���|�K�lh�`����FF���|��26��L˛���'�$P���CRrZ���5�<$��l����^
� >j������
�@FMV�������f##����oU}�?c��˪w��о�A�s鐮4�����BI����F@+��T�z	1Q�>�U��o���z֒����Q߬�iC6�m��(NvT�� ��U����ɴ9�����H�k��W�I��^���8,��m��}X0��F�MNB� &=-�����d�󬏪�yϛ�5����������
NQg��ɰja�`���:��f��,f�̀!�Q�-�q)�'fJ�4o��	�-[���Yb�O �T}o/ i���Ч2���ÞH ��^�o�f5��� ^B̩dҧ�w�^Ǯ��������
��`���!B_B����.x?_��Ĺ��_�'i�_�����Ʃ
v?��]����������q�o3|H��P��2$�|��[kl�iQ9�,�������&J�@U��w̌�Nn��un�-����[<�����x��^'8�����I6��"��V������`6$��0�������G����U��3Q��x&�}B����ǂ�� JbXV=)�i�/F�[��8��7#�cF[e�==@iՁ����u�/z��M�6�PH C�C��p��~{�g�n�`C*�s���$5����͕�`��T�M�wm��Kv���)B��٦ |�$ގŮ�"�S��N&[�:�?_驺g���H��
rssf�YL�ͧhYA&{��+aǊ7�������e��-? ���M!����"�r{f��A�������r�	�"���6CZW�o�7f�!�Owf�)/hz�gQ(�r��{;	@����}Q��8�)-+C �5�*��z��iK E~>(8R�r��3�'����|��M�6�T@���1m2���R��.Z^"*����N��IT���y
*e�\����K2�u������/�4�*�����j|�}M��n��6��Y1T
ȯFR��	~y�a�x+��裢/��biUl?�E��������)�uo[�����Gm"�˟M��O,VV��;z�؏�b?���&�l��^�'
�'{\>�6�f�H8��&�}������F$-�,�	ȏ�����]�S��;�Q�,�.����� bLj�&�۽���L���1"���T���2��0���.���TS���s
��;8���sC��4G]���L�[����ҭ%?�խ�ݩ�h`(
��w>�f��	��TÓ��[ǭ���'{��8��dP�55��C���<���� ����U�Rs¬�ͻ��/FEBI�r�_����P�~�H[#�*&�y��^�{H��6 ~{�{�%�s:V
xN.���߭�X-g�醍N��iܪ�g�T㕁�;��h��xG ��[�UW.}H���߁ر�IϳۢӾ�������ls���V������"�Ņ;&�+OƏZ�o�I/��<�ř��G�r�j)�S�GP~��d��~f֋߂�~c� x|~yy?=�ݭ���-,(�����	�3�2���KVD���.J�����Ӓ����V�l�;�H��1�Y"
+��Yj��OX���uu�B���b�t�����!ֿ[/��Ҟղ=�'�3�>9�0�$�pf�P~_u�T�����񛚇c�N����9��<mQ}��1E�&�V���uboM��gk�-*kg����MQ�� x\sPfq%��ۦg�,L`f�V$g�&�ܴ$��cg�KcQ辪ݒ�C�����}��<�0M�@����v�F�-W&��sc�A�M�����vo���4�@�S"���ʝ�����۟Ar k�2�`?%��.����Y\f�mDLazd~�َ�w��hF���F<�]�)�O͡������Q�Qp�Ic��wnY�w�W#���gC~ȟb$������4݄�0=T2��f��:gb]�h���_h�/yJx�1}�ʹV�(\��7i׾���ѥ����/-/))iW1[*)�4:���Sĵ��ig���N⓸����������}��G&"�+s(Sq��:���`�����]5q,֥���B�i+ݟ�~���)�߮�M"�koW�t��dsT�KF �	�lc���w�"A�����ˏ1��}�Ɇ��z�-��h�!�Ϗ�"���y����A��H�ڏ&gC������F�v�n/�5��W�69.�ǯ�oQY�.B�[q\?�P+d6�)굿����-�;���v��bs1���'X��-�<�,v�������)�g�Y�H�Q����4�B����蝧���6=��O���}��?�O~�a2�WPX&��'C^�S�b����VU�ʏ�+�"yg������2�K�Yg�z
:aP�"����_m?ا2b�r�'(�R���*�f�r'�f>[HPP�X�Ր�����qR�������r��J�Np  �O�#�B2�AQC�S�����P�ϖ[��s��URҜ&x>���}b�gsl�'r�7�y�Ec�IM4*wt����p���kE�G����"y��\B۹60?XK'��t�H�����ة��B,"���	�^�dcB۴U�Gh�+Iw����,������g���l4���a���MQU��-���Q��f�_�~�)�0�䵴�]<؆�g�ZRߎPK��Þf�4u ���Y�\z t��(�g����c	�91e;�x8j����ڭ���.?`[\�(=J��rRy ��q�^j��F*Δ�@J$��rՙ�+�
�Z��ׂ(ORH���-q��+��w:�l�D���D�~���층���0�`]�J�i�VG6�Y�Q�}#[ku��FR���wT|yy�e���A���=>��=tc���[-����~����˦�"5�����G����T��)ξ~~�W�*�ff����aJ+6�����:%�:%_?��z����=oiKPT�M�����o��XN�˓�A5<�u�Jj����E���,''7���}��}f!y��Ԟ���K�'�O23��1��?\�/���Zj��kp�ڥ�b��r�PJ/���p���ۗ,����#	=�f��d����^���!�����-S��j���O�@����>����s9��%�kF֚�f�L����[�d�PlE(���v=t���B� �����i{��s�0�zEG<郮V�Ov�#�Z�6%�פ�7Cm���1��
�ϩ�?0��/3��T�n��=U��>y'-d׼Y�*Ruj*�A������cM�����b�WɈ�( �$T56q��&'�/d���c
W�uzcO��Ч�K���Upb�ׯL�ϹȠw,,���\�5֐Xܠh�&Ƨg�В#�77�D&�9����_ۯ�
���1�{^���e�T�B�o,C���빼�#]Mc����D��"EϮ�~�6�vXPN��
� �����OGp<�����*X���(�r�\��,��¨�s_�����R����k땯���ŗ�KKK�����U��V�����C�M�66�w�?�u���z<�e�{�-b�w��G�uuq����匎��g+Lͼg7��I���A�%�1��	b����2q^n���T.��R3���K�-ǎ�����L]ZZ��:��?���=$@s��!�pe��kcG�]D?���1���6��9�˝��������I����ЫgILc�h=�A�>����1n� ���h˵g_qZf���/��F<��M�>*Z��eq�3)`ڝ�M�@���ƹ����:���;��|?���[R��Å�e�����,x-N���'��k��Q�M;�i�gҧ�>a�HABB�����]�Ԕ�뗠�guC)J�;?�X	G���/ܜ�<��d�+��:Y�R�z�6����p��������4E:%\��x��  f��s�gk��;z� C�*#.��/�]Er1kBi��!�o�&��[���ʅ�I�k�Z�x�̃a~��	���a�2�d�,�Mj�b7�����d�@��O	�����e �F"���V1\��=N��o�bz�E�/�J��{��D$ͧ;ס�/�Q*ϞˋF:î�n�.�b��c���*�������/΋�D�T�%.�uי�[^� \�w�4�q�+/�i���`f��/�49��Na�D�!5��b�&<���,�mHe~m)̀��ڿ�½3����'�wƖe {e˅��ݹ�G�FMԀ�{�7��	ikV��*G���j���b���SE8��e�>�A�uK��5�4Z>m{HϠ ��4�Wċ�5����	9�J�`+�����P��B=�0867���N�[�P�^�
vo��3f�L�5]%i��)���m>^HT4��p����47w��@��C5^?P�^��ş㶢:|c�3�O'M²[?-���g��o}}}	ZE��9��NP�dSII	�Q:�ysl�p�h�H����$����BM05(J�FT�319L�"��Q��>^U:���	N֐q�0e��ƚ�6�E��K/�:�a�xF��@R���3̝��a�X���H��'����L�s�=��⦸IE51)�.��p���ƷC����<��q�E+�eJ+���p�}y i��=�M�.��uN�3�9�r9?�?��rT��SЩU�"Z頳(;�F�*\�j��<߸�=���q�|w~�G~s��8��5ݿs��1Y��㞄dǑ]�6i8M�E�?��2��ňw��v�4�9�S�9�>���)H j+�"�GMO��Y�0�`�h����~�^;ȏ�ZWz��M�Ǿ�Lj�^��(뾤��Ѭ��*G��	�L����m��#t������+Td���Y�Y8�8V��ER�`lQI�4�g�7��!6C�f�o�j@�Xח���
���W��b��XϓO�`G0�b�t�a��e�.DMٳAĜr�+++�'�8�
����O�%�h N�:�F�?IO�%OP�b��j�
ʪ�x?;*���I�j��� ��W�D2���Kdzy4���!�)��IŬq���1�r���� kq���,f�љp���u{۟)Y>����oB����{B��^��[ �A�w��v==�o���ill��*���H-�W�@���8[� �]���F&�r������#�2�+<�S��_�4�Fv���4`�6�t
�j!��9���#�{��_��+a��.��X.�~ᴸ*�������3ҩ�e�pi��=�,�x��B��ژA�ej��2N�_i�(��R��M��1P��㸉��r�=�r��� ���ݮgn�M�YJY�6*d�mK��[��'���;Y��4?�����<��LK:�s@g��il('?�*.¦���6���7kw�BJ��Y�����݆͔gw44�M�0�&R?55�>���p��6�dQP=��e�g��%�&E&7WCX__���O�%UU��L�΍/�FZ�*���?�����W�@�g��t0�ǭϷG�x"��l��.+ߘ��G�ES��(�;ȝ^<����LO���'*�~�Y[����%x<kb���ic�՗��c�fy:dmL�.��)��x�b͕�߿���o��:~�B�z��3��%�_0�'(D��)�
6b<u�Zm�)��,ە��nk[/�9�c�[4��E��i��JOX������s���5���ڤ�4�Q��� � |X\�no!1�s^�C�w���'-�C��k�>�l������pձ��m��R��~b`<����Xud͵��W�i0���L��5Ng����5�E=?�h�V�5�ޱC��W/�,�~7��$�U~\ss>��$QO�|1*�x��2�JD�J2����]�XW���}�͔�'dz���Q��g�Ⓠ���]�fл+JyK���N�&�c�b{?s��\L����w�s�^H��I���p�T��������V�~(��խM���s�4����m�`�y-���P������^#�[/��m �%矁�=2l�lp���'-y�x���w���]/�Fm��w�% ,N�;�Ⱥ�ե�'>����>�=�z���߶�xk]������s�����(K#�H�Ji/uj&u��]�P�dEW0&�ߙ��B�pz'��|7���?��U%Z!:��Ѭ*q�:ؽ/J03�_"��
Z��Y�2��<iA��)&��ڛ��iO����o�,R�q�t�cv"X'��ɴP�py�����I{��g5U/�elT�2<�b2��������0��ppC���v�t4+«���LsG�FU�.�A��q��*kj>���M����3 �F��#ej/TU�[=���z��e�N%���G������RS�DZ g�7a��{!|��p�R�޺�	� ƽi����1���}{[��&�$���pJ��B���C2FG�M�F\��.<��6�rlR�P����\ �����6-�~��VQ�'��O��&�0�,R��Y$�.� ��Q�����	|Y�Ђ5/�x�YB#,���q�MD��Gإ5�t�+}���P���i�������ƕ�uz ��q)
�o{���5�c��qf�n�TgQ�4k+� ��׍��Я"�w�ъ�[�iŤmt��ۅ��B����	tQ�y��!��g� N�U��EY׈� 4qȩ�_�Q��;�ׯ��y���'��ǫ�X�Ť�]�p�;��K&I�;N��ޮ��ωK��o߅�H̶�9��ɛ�F���D�oW]^�O��TEj��,C�?	֌��z�t{��F^6@u��b�jH�H�-���~�pK
����
=6&r{,&�i�X��tꦌ��5l[�,�U�9������v�, �l��K�B;ś1�u�l���MgVzU��W�"x�o����Svе��,�����ͽ�{��&p����2U�C���XO��A�������چQBR��Q��NA�Aah��SJ�N钆A:��.)��n���������pf]�>c���M�5�*Ua�~�p��2#�wJ6��1��,:1�$����
����j�i�}ϣ�A{�n8!��x�J�ۿC���)�CTXXX�v(QktD����腩l~�}�����d�d�Q�:���U
��?���\��e��74��kqc���DFm��a�~��A��",�
P�b�p����/,��k
��\��ٮ- ˲��|�.���2��sV9��|�(�Ӌz�nd�Z�ۤO�c#}/��'���^������f"m���hd��V��s C�}C���sD��)�$<�=�>l�7��(�1~�8~�ȝ��\���ƀˠ�ͫ?q������S�z� tt�!B��2���&Y��Z�������z������G�#F�E,�3n�xe)�w�Yۄ �)��]�B
(LC�����L����I��e��F�+�'�xiv����OmZ��C]����`�v�G�\_v��a�y)��{~O��H�	F^��KS���/]G�l3ª M��%�^���ῥ�n_�Ev���pw�?T���N1�2HǨWR�gv��z�A2��W�bM�$j�~����n��n>�b]�`�a@~��`o���l^ e|a�?D ��Y��1�`��N�8�n� �o��/1v>�Q��.� �>�_�?D�rQ��H;�cK���i*x��G�C�O��7$����j�����6
��(?��\ ���bo�&+"� lD�G��\���֣f��;Q�N��v+H��ijc���$��K��S<;D�>V�����R^�Ƥ ���5��(�p	�����(��ܕS����,6}k������?1%�9��j:�t`2��h���!×��:vuۚ�E��Nc^#q��P����Q#����;��B�_}cn.B��V}��A�
�%�77�l��Ǒ��|��.߾���"����������>-�ã:}�#��x����HrWG�B322�N@	�^�H�\.9��\I�^%~	�0-T�(l����d����8�?�KlőD���[��d��ϼ� ��������Y]�}6���O���D��u3i�`_�j�vM�?)�HHͣ5ƿ�,+32(���3p_��ӊ��V�O�%�+����ܡ������ I^	�(@+�%�;K�K#~�}����9Gʧ\�b5������-eaX��^J�wP���9�鮀=ےW����S��~q�/���킼�CAV�^w$����Mwg\�:��g����'�i�]}��#?m�s��']�N^:Bۘ�5.�w=�7�� U��X�������"|�QbW�.�׼���wp��4<<�1����I���&�
?7�"����U"�U�t��́�p|bj:T��A<)Sx�Y��c/�4��Y�.]屫Ӹ㵐��G�X�s�]5��'�`����wz��},��n�|)#D#��J�%�ġ�X���������>R�W�N�Y^!ۭ�U�b�z��H*��s}�O��i��[^����k����s2r����p���*U6d�����g��ݎ�_�W;6̴,�J��h�zNj��y���&>����`�u���!wiZ����f�߳1�i��اy�\��4����))K�����:	�K���kR.�@�>�����js���K>����x�JD�"���R�����M"����!u!�����^� #�����l��2���Kp�Q��mX��;)��xn{:�����Z�%W�B�	<�����}��?�1<O뚂�bk�&p�@���/��eCJ#�]*��<�A��p�P���Р�!��ɰŕY��M*K0�W"��7#c2:�l��ڬ�6�}C�OX���^�.'��ه\��5:��CbJ9)L*|}}b��h�C���j�N�R,����y�^���e��ʆ�c��k�9�X	 M|g��
nu���y�����A�?l�Q�^��\Y2u������=6��ʑXܑE������vw}3[G���U���\�ZR\�9�j��Ď��_����`v�do�h�NV��:P\\R�Yri��~�V8,�Xh�7H�T/�w���د��(l)a�h�Q�s!:k�-�fe�A��yV��
�B�))����9� s���H&Qթ��3M��g�B��/�R���Xt������!�j�d"��	�N2S|b{<����&{c\j*3���ij8@���	�A��TP��r��$���Ez7w�N��+�6�9+�TP�7`�x���ޅ�U�#uvv6�R��U�^���ڲ�aV���q�������O�L�
����&����Y��;dz�����O�(&��Imgn��Nt�C	q;Ġ���xmt;70�ۖ�D|�)�|�d+�;��c�75mk����[[X	���с<in|!S�k��;{�}�|k��h�aq��\�PrU����Q#BG3��3Mʞ�"2p�J�j��L�%OS�uJ�c����vb�E}8�:����4G��22н�I8i7���R�57GS-V퇅�C5����+�Lcޝ1���jG������海Eb�^���|��(�*�Qu��E?+c���y�u>Ͱ���ߐ�ޒv��sVF��E);�v��*���.���p>H^7l����t/+!zD�G�l}���Q�2>
��a�cz�oKf�-���N޶��׽j���.��z�����a����m�or�\��LyB�VP!��ۿnF%Ir�/�����;���C2%.���\s�ejCq�޳9�j�3����-��B8;`y/�>��6�M�T���������蠹{I�+}����J�CԊd::�KS�,r�WQm��lgY�k�;h(7\�}�ޏ*�3j�M���8�8���$�i���,:j��Y;<j�2K�KB�"?8��xHR.�,�(���yO,�h�+�����g=}*E��\�rA �	���_j/�Ş����QS�j�5b�]���4��/}7��>V�p_s��D���2��4�@}!I|� �Q#ǱUR��_]g��=�E�&.�v��$�=�׷�������.�il|e��y	�b.����u�D�N��9��x�6vϯ�4���rrr�RR��N��c��T༛@>��0?S�>܈'�)���p���V��̜5���:��켏K��
�"mU�Ǒs�avz��f���=��=?�낣W���6$�E�孛ە�K�ҳ&�N��z�\�&�.�:���}��T��)��-�iN����#�|A����k�N+Z��3���ǰ���;.S���G�8��$����q�6<��L�[����p�t2�>��|rQQ�S77�)g����T��c����4K�ٔP�	4��4L�as�+#�@�К���r+����7�D| 5����6]�r�SZ��)�M�l<=u���68��6ihZ���[�:x�O��ZB.a>�Ɍ!x�ū�UF�?�Wχ+Y�z|q'.�u<(z�्MJJ*�v)�n[辤�xȬVX002��ly5�w�u �,j���'ʴ��I���� ��_<��^��&�sY8&�K6�S
����ċ���l��I8m-�$*�n�!�@��-���
L�����"�_�fM������P���.�/��D�AP�E8�);e���!D��5�9�n����7�Qÿ��F��8A��\w��k��Ri��#����Ś��)[�B�T+Q\&Sab+壼��e��ι�n���w�B���v��s�ۿv+}����?Џ@,�WF��}3�b<��ϛlq����6��8��g�$��Qj�h2r��Q�Y�P!�BXճ" j%�XG��8*�� r�̂[���j8����}��W��P�{�P��ޖ2`�A�7��L<�o���I�,��w�aN7a�v�7�˝=g���(Uݶ�����y=ޤ�7h(y�MF�$�Fx�Q7�z0q�Cq$��5�w�&��4<�J������]�b��3�#�]i�ۡ���Ն�G�/`������(��3Ieī���<���^��q��h�\ӭ��/���+����_{}��2��)��}C��E��ݍ��0_Z�a�4��y�\Y�X����L�N�UTT����V�'rx�Ƽ�O��!u�	�<�
B%Ǘ���>�kǒzt�� ʧ��IbX;`NZ �ą��MɅ{����2-�GU��g>��ʒ#�(�]Y}�.����L�%$sPS
�|p�ԐD� �M�e���/���ĂJⳀ;S'�>�9�� �P��}���ǵsm� 'ܕ/�+%��3�+۔41jy�O-�7$e�N����y���%�E�S�g���C�	�����@3tA�}��͍6͞�|����A�~$F���(:T�d�e�L|��M����	m��i�^��?��ݹSGQ�!S��g3�:������X���.hO�o�p�[c1سu����WL\�8Yʢ���b�?�	ND�Ql>�:jX��
q��?���%����#�W)���W^�i�w�P�WZ
�d�5���J|�ŭ�QB�� .~8	���A���6��D�M�Zc�ޔ�Lx�vґ�6S�&�_0F�+1d4�q����,�	u�P��}��� ��5-M�6m�7Lk��1%,b�w�'���3���zF�^��L���&V?��ץ�ｦ����=4��m��N���I�����g�������ܐ��UF8z�-���V�E�Xi�	IU[��M��;;�5F��۞��QĶ���ok}��������.�b{�,9����{�v���,�%�Dh�^��ib����CӸ�3������$ciy�6���P*����O��t�[\��������<(���D��m������h�ֹvy ���<�Se�594�4X���C�Dͤ���,�)HT���Iw���}`5Q�?�=B�U	j|�/f���^��q�A�Sl��p7+�_�4;-id٬)G�
"}�A+<{� ~��as^�������8��ͅo��6ܦ�c��G��BW��7�}�J�_J��8o�+ ��,��r0[.P�t��Γ���v�J��(�S��PoZ��"�F�Ϟ��\-�w5��E���F�C�� �':��A������W+&�i����F�bO7L3���*����i��,����>�޽�s��UZ��I�n��[j�ZS�CU�H�	nR�����(X�/��X�k�f!��j��m}R{~�Ph����2�,ږ�!��PvU�*�OG�*Q1l��s�N+�I�������r�$g\h�sYVq�?�@qb�aA�D��ʝcn�|�f�W[�gV$$!]������V�{�Uqw�����]���w�!�c� ����p}�Zlw��锠\� ,hN��4Zt���V�n�'�W�}�	�U�-j����o�t9�1!3X@�
#a��1ٖ�;]�Š�b,�u��z�/�Ď�fA�?~���˽�O_�9f/"�0!zC�C�����j�X�`��O��ڇ��u�,w�]2���j�a�����<:��Yu�ygNa����),���FcxW���{+����jl^�xk�2��ޚ���@�U�umi5
E�gQ>�K���uH4:̯}�-�>�S�m��r���@E���C�zuj�:q�\܉MLA·�9�j��\�=1)���V�
"��<��«K=������L�g#��10��ph9'�.F(�@u4 Fh��Ghhe?Q6��<�����y8�T�5�`�o�|�/Rd�������hz����{������o�+?�a��RBF� �$�k����j%�w�"?�� J4)w���ͥ������g8��l��k�S
'� ��^���W����}O�'��~X7a.5����������脓(��P�Hdhoω�_.�7!0�D�w�jWB��kB���F�ӱ)�����xyq�Ț��<~�Jo��
��	�8G��<�9��oT���7�����:�YC~SD� �����B����m������Lۘ�_�x�@u���Ńm,�˻���!��s��LV����j�c�o��P�cC��`����W�V���n�y�����@��ނ�8%�Q��l�U��j�E�Ǜ�	á�i7�2k//��p������7Y������^��iȲy��Џ��t��:U���}����H(�n=n¿ ���]S�:�%��0>4�/���7i�Wx�TR��뭾�x��K�"���f#
v��_3<Ű������H�!)s���Y\Z���dڀ�|x��y쐼?zz�b�%e[���0�ipg=�����W|�:)魤��M�vl{&5�֡�G�*ax��&�(p�ٓܨ��6��-��/O����N�e��x ���vJ	��{�5���q���"d�æ�mh����k���}�G�������uE5+�Ϯ@N��ЙF�?�8���SA2�X��ɘ6�|�7�Z��!6���g��j~:~f�޸>׵�j�FΏ_�Gӵ�6�r�@<������b��\׾�������R��" P���8<'.���0yC[<��:n�B�/��O�zc�1f;\E�aq�|DrP���j��*DϏ�s��.#L�~DF�;�+]�����j��פd� �3n�ՅøLos?l5�C��5���hnM  ��-�t�oG�x4פ���=^PR=��H�/S�3z�!��*�޴�����;#-�A����^���Ō����\|��¤����`�P��`0�ө�����~�@��3�I#��<�7'��jAɹ��a�d�]z`��� �+a�و���OC�#���vy��fV,w�e�%(i����&*���rz��:C�h'�12r傿�{@�����XJ�~�Vd�h��4#�j��iW�s`VCN[H�K�{<��\��Q��TfV��]�m^��όc��lF�!�9ل NF�5��ԧU��~/Q��������ʱҴ�.��|Rz���5z1�k�����'Y�7o�"�R=�����|_�4��^�+�!i2\��I�����p.9fW�&ط����DOb>��ǓXq�zzH�&��	4x�d������1e�K@M<�E�p�x2utgw�;Ԕ��/�x�5���Cq�{q��`6%^�(�2̜.[���t�ƴ��էO�+��,ر"�b��U����fy������6E�O�����[�9�8����~��}!)��$�M~���hnc�q�v�L4�����p����q�D����Nh�1Ud`ꯧ[py��6Z�� s���m�J������=�����>����6�ΛՃxOˎ�t�+������ҫ�#��ڠ�Ј��w��x<d�DHn��i��g��o+g��m9b���nm���4�����Q,�iba�\�SV	寰��Jb���0���e�zx�+����"8"�M7�5�����s�W6C˽���%P��Ύ��|�9ʸ�����T/����E��=��`�6Ϭ9�
�8 {`��_dAA��Ke���;F��,Ow˅ee�lӯ���I�{v�fFSK+�ʁx�d`�z��}�LM��~�So}���]�l�\�p��C�gW��?�_m�0�}�y舌~�pZ�@������^�^����T�4C�:[P�e�ih��M���݁f�M�ZZ&��X�k]wdQ;����d��4Ѣ��}�͝�ͷF@N���������J�u�l``g҉�ߥ��Pbv������z�� Ը�Y^��Ϋ+��_=���~|{žv�3N�C+�Fڂ�����Q���Ғ��"̎��-n���9�|x���|��H������3x��n�-��*�����T���i���_��D-��w���{5F�=4�4��ض���kT���������Y�6-fU5��9��ן�=o��d�u�4F�!Л~�kH���O����m>�p��-8+��\dl/ʔ�J�~�o/���CԟZm�s�_<�1��0��yZEM^��:�c? �����K�I!�u��#���LRix)��qI��*x��j�T���O^������ȏ���)��u�~u�i����v�d�f[zQ0���q3��v傄"�d��Y��<.���qR�|A[F^7b�?~�D���{�l.7e����t~�?[=�H�O�)�.��,���r?8��^t�p?��;V�{/�4s!`BѰ�j���V"�U��GbQ���k�%o�Y���B�}%a�O7q��Y38�ٗ�qv	\�v������f0�{���ЋY���<�D�b�>GJ�6�������������S<�F*�"��ݝh_�-�x���x����a�5�h��"��`n�Mr�'�MV�c/���^��@��)�6 {Xx��^I�On=6ru���;lY�l}� \�)y����K����<w���)�s�ۘ�-�������}�A�yۢ/���ꂮT�p��x�9�L��@wJ ��d��}�)#n��4�ڃS��=�:�X����r���k����ύ뎁aa�BKo`�~������7d���:eDj=ss�L۲S��BQ��-n�ku㒙��^�s�]�c&�E^W!)S퀽�y�s�5&�'�""w�Ko0��*�$ܑ?���lʴ���mtd���j�Kf��p1���Z}_i�M\Je�w]XX�=�7�J�R��)2I7r��&�;k���H���h�x�'��i~D�[Z�j!����B��F�[� �D�w��e	�'��(�e�jO��6*��+���N��8 Q�&�a��&Ҧ��{ۣ�;��p�u������ԷX�����v������G(�n\�݇��C���k�ϓ��=J�.J�Z��2���d�.bS�b�'����춱��3���k{�v��}ԶY$�$EJc�K7/����N��I�Gu�?���#���R�%
edj�u���㪓��>��ڥmo`���[�ι�B�o����Fq\���T�z�p�t ���Ti�&�7o�u��䄅�9�\[��]���e�ˇ��o��q��nH2�ݎ��܅��f�b��I��C$:�6=!)z�9�s�d��?�܆�W�ܤh%�|����R�Ϳ�.%�R[ØU�����yf�0j������e��j�a�"؋{��}��,膂�` y3���n}m��<����{T�@K�ׯ�5�tb��r��yJ@B^f(1/���B?�Z
�w�V_{r$a׵״ԕ�i�|������a>���Vg�OKN.��G���=%���.>>���J~���ᡴ�Lkk�x0�_AU83�l�O���f���Y]�PXQ��^w~�|@#>^N��#l�����s����3���\L�T+�Hw��z���?���?
�!*���.V����z~d�Sc��9��oOM!�ܬL����vK�P�~Ů�4ZW2�H��jE[ß#虀��ݷ_�T��^H{�l`����k.��_-��"�����|�|y�����<1e�jz`Of�ɮ��,�ͻ	����zv0pߒ6E?��?�P�*���~����~xk����h0�0h ]�s�}��s��ޒ#W�cJ�I���#X��g���R���X�����2Q�
?3�;��pw�#}4&�&3>����sa33���}�"��������Ea2���Uo����l|�Ƃ.��jĊ�@�vG*Ed�os�9�څ�l����d�^p ���g��B���m%o���LZ"�R��u�W~!9�����=����v�Ff�1�So�i7��+�0��6��k����d�W�_*A�i0��O��Nv4羿'm�Ub-\D�Ծ����K�mZy��/ ,�_Td��bj�fxb ��B���^1���Q�h���-XL�%7�)�1��i�������8�l���OOh�\{ ��Sw���ysǀ����Q����gZ^�{��xMT<�<	�-6��'I�;X<��~��\�TY�Mg��Yͨ�J�%�l� �p���$�����)�o������]��D��eK(l���)�&���I���o�L�z}}���	1	��'*�;v��Cܾ��P&�,�9���8�8?}��+U��MF����H��3/�~��f|�&�X�lB@f{�;���;�G�A X��~A����m�).�Źs1:�_c����������ak�ɽ���[�r�\�H�O�}�8�k����ST�a�t�G/]���ĕX�~V�&@g&e��C,�Ȉ�{�Ģ+-Z�|��:W�SW�A?Y�w�J%u����r�G;>��{I�s&8j���jK��&q����ή@��6v�f6f���i|u�mykF�,<(ê�]�4��?�o� ��G�}���gW�Y�I����d.N��:7��:낈�%��`���Q��e%���Tt	.m�z0�Ƃ��ʸ��]旴��G�BJ�I^�����<�޲��mص2-	@?�+��� ���|�{2�|u�>)&
M�`���g�:L}k����-�#�f����k�O�r<�H-��7�Ğ� lU)������TQ
8%�z�x��t�gR���{��}r�4�+KĔ��k�7�$Q�/>�Қ��9W�告����~�UC�	{$��L�%=��ߙ��.��M��Գ���Q����U�@ݙ;:����a���T���B=���n�����.K���[{��nb��Ζ8�� /5�7�8g'��_Zc�L��.#X.6$��XV�Gɽ����?['U�
n:̫.1���q�(q�ynz���Tc�����!���R�ѯ4��	w��:�P�L�:w�(<�U��\!��/�R���P K�G���!an��C�XCJv�I���k���E~e9���B/uǸ��yM?��L�	pq�\Z�aJs�u-C��j�N�1�C��b�M�6K.�Ő�O���Zc�5l�)�T�œ;]��P�D{�y�y5�2w�W�Az��گ��pF/ʜ�X����@����E��u2X~�}ł���h7����IfM��7��<�/G��6$�
E����<y�~��%�׹g�<��/&���#���X�i�!Z�BJ �Ęť��߰�r)�-�뿅t>`Gↁֻ���1^ab�����K�	���|l,���7tŸb�k3؋�F����س4��G���=<�'�OK��ūR��Ox��rP���ǝr�g�{��;<m�k�����ȶg߾"jG29/Қ�I7a�r1b�ݜ����ZN�Ҫ��ޓ��\vm����),��nR�/q@qd��4H�	�f'�z�'F\���TX�q�2oy�����JZA!�
����ի�H���W����/��r�'J+���C��RcH(�u�K[<e!ca��e۞����ãǱFsΗ�-�Ce����q��+��p����5��u��u�8�w��l�����o:d�_�<��y����4�W5p%*3�\�7聍�w/�|�g�άύ��xq}}�����N@'Ͱ- �8zaƓ?�����~Hn,5���!XcY��aW˸H��-���b:15,wŭsE�}|?�),'�*v�w��	K�����Ǖ�l���T$��dq�2�~�VV��ONK_''��uz�X_�*:����a�m!?#�z�q3���5���G��q��k��6�Ć���I1��O��$��G�`Ii�?3P�����_mX��&���F�?�bG{����"u��N��@r��q�!h��������f�r��G,< �=�g��ma�3�a�B�;�J$�z�^������\��=Kr/x���>a ����xo�}��*^��٭'���ڔ(��G2���"����&0}�a�i���x�4�[�3�f���_�7w+�P�>x[S=y�
�7�گ<�!˃�i�n����F��$\0%�&%2����ª܂ZG���g�$��p%��cVI5{ ��+g�1m���#
�O3pYUFXW�Ͼ�=�X��4���{�чxZ�ƒ�hƭzh�I�es�&�l����ݠW���^�N�2J��)Lw�+��K��r������_�]�W�`�;O���-�3U��~4��X��b�M�f���bm��BR�<�[9g�L��r�/˂������MQ���r4�ť����J�}k���o/����õ�vi��?	�� �2C<t��a�j&��~Á��-�d�kݗ!E�<􄆪��d9m������+*�:��V>�����Y�Щ�Tϑ��9hd�7@q-��7Y/��_-�Xr�Z��]:,GFb��b��oS�\r�Vf��v��p�x(��c�r����JC�o��/9Efݻ�������yy��#���7������^o��L�w'�O��"�T���*�G����
�C�'��F��B�b,j�|:�#N]3#�ĵ����=��ψmӯ6��\��X�kt�I�9�~���(5�N7a?{9DuЗ�lX�TY0&��	~��Ux��ֽ7&�0C6�UY��Wܼ��6O[#dd�����	�rZ(_7k�ÝD�;n;���K)��B ��6�[=Eg�h��	��3Ew�o�o�Q$�d�#��v��g���/�����B��̀��z"���d*����5��r�O���Ar��>�h��n�����+znY��[LJ䕺x�*�/��HW�!M+;C��w��y"��@vl9�+�Z�]t���,��:�i�t�T��%hT�ц����<޻t�T0Y
�H�-��\�8�$I/��j�l1K�����'�.�8�8D1>���޳��~>�`hb��;�'�៉w*���Q�30:�#�P���
��p5�Θ�/]0��p�:C`M�����2���v	��ω}����)U��nR�Q�&����T}2Q�ր�X�%�� A����k:O9F�[�d��$�-�u������7x�a�O���l��t���	����E��'��}p>�+�SA�-Q	���:�Q��{���gn[�OD9e�4�@N�-��7����l�r&���݃��q�_�����Nm5���)QzR�z���q��v����%��Ǖkq�Ŗ���u�����Y�Ý���mW;8|�Uk�r?`J/����t�5�!��9�A��=R���jϾ�8�c�ӗ�;s~p:��V�M+;[�����Q�4�5�>�͑�d�ؘ�����BLOW�a�z����r�eѣ�a�����;�B���/�_Ƴ8���|��K�`�a�p+��C5�D�n,9ԋV�����6"E7� �� �|W�e8c��\�F��-�Q��T��&,4ڗ���F�n2׶�w���Dqd��cߺܟ��u�L��90S�w0_׮���e`ް?c>_�2��$��FL�ۺ���I4����a�/���{}UB���$�.\�B�B�vm.4b�nUd7�A�w����In^���p�c�4/#&����LLM�s�*��+m�0VQݡ�b�l�{�y#p�����U&kN���Z.[��+h�&��P�KK �Bհ|��[`�r_�[^>� ��13[\�G�����3�5�qB��������^�x�|���0��z�98�X:�RE�,0b0t�����+;<^ݞ������Q�%mW�A���=�a�+��&ey�T�pL��uj�m�t�]����`F �������ʠ-�_-AE����I���!��ꝫG��k���َ�%p5��9��6��'
��{8��{u�����)�^�TNӰ��Y�݋��:	1�ޚ*9~\��8�8)Ҹԓx*��ah&T20xv��o��l.�ײr�����`od8�����ug~75a5a�~��^5[�#h���Vk�C�p������8M����ұ���`c����z-"��-�)+b��Q��H�	py��A�ok�:6_B�8],>�l�<W���Z�5}��7n�u�(��**�Y�S
�̚��sܗ�G^B�}CVL��&@f:I�Š�#�� �w����Q_��P-�-�D�v>��Bι�h�vx��FZ´v��J���w��9����!q�N1����d�ɖm�6��{l���}������/����^n�Q}�4�����+�M���ye%^|8I��	[��.J˳C5����fdD|Ik���dTdJ�J�E��~c�g�$�rHZ|I=O�@%���ճ��`����d�u={���Õ���k:K���w<7G]��FK�Xx�L�b#w^iLJMH���G,�x�(�/��3���jLC`�Tv�ElAS=K,XA%me�۩w[�ɇ󉊮�/�Y�ŦG��%�yg��@�������vP��ᡗ"�i��Ɩ�f�Y�! �u�Yd;ē� �;�]py��~UN�]�F�n���MM"H$�@�C��|��L��
'�}4��V�������ʯmeQ�7,x$���kYٝ_�J�%,�(yI���|�Da��;�x�G���Y;�$~"�. \��7�#�=��J�'�]㧷���G�ͦ�q7��R�O�n��|j���C�ƣE�dq�\���'�������O.�rum�I���첞��T���"�Ăr��H�$rթ��Y�!����I��V$2
���G��T�YOʸE��w`��h�=X�-��հ��Ų7����ql��0�T(s��q%#���>����[\�M{����>��Q�6��<Ii	p��7&
��[nh\c
[nk�����^!�~��s��J�MN���� �!�&����R���u���	��T�_8=�:^�\����i�a�S�=�MG�N�����ݫ�w����Y�M��<�vO�x���}=�������!�*6*
��g'ڰ�����$�ʶ�sz�}���_��	���(�J�._�ז��~+vCn�z��_�D��Bj�2|+rA]�ƃ�Z�r�N@�>OaG��H����`F�'D�cV��zv\6T��E���t�ms~F�t�=DI9x�ۘ�Y;��1�l�vh���l���D�:�#su�D���,������Z�*�	���X�e�T��l����'����ԑnCp��U�~��WF�_��6ˌ->&�M��/[�,pi*--�U���Ը	L��\lm0=��t(�Դ>L�b�Ӹ��&){�O����6u�>X�SXޔ��������?�S8�tf�S<e��������@�3�ג?)�ѝ��o6	=y����x�'�����ϧk|���'���C"��##;��qSMyyy��1W��6�e�Sl�6�1|׬c.*���:����-�D,�t��> .�����S���'��5̜]���d��x���c�u5���+��Ë��EI��~n&k�X�k/~��Q9�6�3�F���M��T{���ԤGC�]�^Z�r�;~�Rܣ�ǐ���_7�aċ�X�j��S7na�Mvwy�w|�s�>�[�����Ebff�����őL�&)�շ5� ��f�<h	��,&`��Y9��=���x~y��-�y��^F�y!J�:���>(7<r*���H��������d0% ��,�pC���P�F/�f��+��a��z_��&pP��U�qY�I�/��������J����c4�93a~�}�Ō;8���;�p�/z�M�&�uч^�������>����{AsːG)�y��۷m��x*�**.{bZ::�#0����q�rL�] _^�_�6�_��ډ���T����ߊ��qb&��g��W��F2��k�#R�h����?��8�E��y�i^�L6�BlA�y�<�}�K�[�Z�ƨ2�'�pE�Y�^탆�	��y��J�?m��ף�OXG��^�F�6C��ֳzEEA!a ��>�J����9��i��PkO�AрU�UT���(#.#�Zw˙��%G4R��y#G01�"n�b�?h3�Jɰ�v;�ִ��=֍�.3�G������i=�x݋v�=>��ݶRv&�2`��g�}⫧]����F�8�J�u;J��$�.��2=-2)�g9V֩u�3����GI����L�o�\�8�u�I��.����\��m��M���g~w��d�E%d��dڀ)�M%����t> �S�l�������@,#
NdŸ���v<�d*�qQ��M#���-k��Wd\��O&�/���<.Z"RW�����F��� �W][��Wx���e$H'�T
�s����#�v%c�pct���=|��`�����Wƃ}'�y>t����,���n��b�o�ESc�d�|�M�z&�oii�Kw�=a%9�Û"~{(����K���(ْ��]{a�G^�ˌ��ͅGhC-��@��ˌ}Ï�`^��^���H�N�O�>���9�l�qC!��~'����"��;:Q�zW�r�ܼ�#�����E����K#b�`D�'Q�����Vx��Шk�Q�N�������H�;�r��4|�a�#pB�xE+�����o�*�<���_���⋷^�������XT�/�;{���R0��D����\�k�T�E,����s���:�L��YƯv���m�8������ѧ(���$+% ��;�CڹSr?��mo�G􄰲�6?�߭Ơʾea�'|���>��[�q#o�+���no�)R��O�~,� 7�A}���ea������o9���3����MO�����bPt��B����}�3�؉Ա��5ރ�9�$���u�CZ֒���e��q�t�=z���}�UQ��/�8j��G�|^�C������7�^d����I��JN7_P! RT���$����$�L��Ҹo��\)K�������6R�y9yK���֗��4�Y�3Q	ɹy�kV�T�eX�[�?L#!��(��t#��ݍt��t#  -�1RCH���R��!�0�������</x�u1{�����Z�0z����D�	0g��S��xTN/��sO���_���%��_mcJԑ���X�N�a��ٲ��HhX2��I��@�) �)}[�AFۭ��kvf.!���Cf��ٮ\��t���ɗޚ gL��&u��Z�q��,\�����mi�B�>��Ij�H-�(�<�rF�Z��aj[�Tڗ�D�S��;�F<F��I���Gp6a�A)NO~oV�����Z�t��Ѳ��>�vP���;!��)}���Ǡ�A��D�cǏ�;��0���%����WrC�����$��X�xM#P���ޑ��m��0�+Y��g�`M�}���-6���H�B��}A���.�)�.�1µ���$�>Z����%e���%���BA�丂^�T����
"�yo��YܢN�<���rÔ&�O��s��{�fS�}F8� �$-&ZD(���M��蝄j+%�w��N�#���I�l���0>���Z��=�(�_s��~ �d��2�C#��sh��?�T+b��_q���Bl�r�I))6�}7�K&��=AZ:	S|�!�6�" ؝lO����V���Nm*�F��P"�����D�xla�naI���Z_2��D��CJf�}�6�/M2={��h+���P��wgdA�jY��{tV������S�\_�ם$�[_Κ�]LⲆ�����ҫ{����Aǫ���Vm�R�{�%
�n��w�w4�������b��wM�L�h�8�g��"M�8�ӠT�	�*�v߹�UZ�<Cn�uy��wa��B�{���Il��т�q���6��Zoy~)������/:ӊ ��w��X���dX(�}�w>?
�Γ xq�����uH*�P$6�B��tR׹�v�*S_�����I�D�>�����R���3��r%�6Ɲ�@�KS���"������ə���-�k�P#<<>p���ycEVX�#>��pk2ʤ��L~�Qo4^�v��� �����ʬbt���²�`)��N�Cx�kvO�lcy��@�k0	�C��Vt�H=v\���CK=�0v�jJ0���k��+��	ӂ��2ؘ�~�D!�n4#��6��;&!\vĈd�!gp��#V(�h�5��0���Hz��'B3�+r�F_��>9������� ��-Δ�W�����ǅ	��N���������	�p�f[��&�T�;�_~�x��;���3j'�������Lac�U�ͼ�}N �+mϏu͖��A����Rm3�B܄*�Ǎe¹�e�o717?�>�_����c����C
@V�K��|D#S�̌��J���3��`��._�W폞-����nX��D���'���\�n��bͻ�?��5�?�[.*h�t��֖-odK�)�%-�:lJ�6��Ĵ���4�g�薪L�I<��}�B�A��s^�Zk�zE�C���0��/~�p�z�V�*��n�S��¬�J�Q�����Ќ��!�p����ö���5�4�%5~F�.ܧ��ݏ���ܰ/�+����ݜuRSU3hi��B�v���ym!~��Cu�X6���'n����6iPϽg,|�E+�WZy9C��f�<��x�0nQģ[;__��Kf�������&��Ć88��&��`�D�6����5�ܰ���Ү�������h�p+������1`��[ʡ��MwY�SK8�G�xKZ��J���	Ji��oC��Xp܀ ���#�2^�t��V��[3Z|m��NҠ�d�(T �z�;���;d����h����שWֵ	0:U�5��o�����KzLo[N/�5F�`棵����E���Gy��y���E�'&����0/�U�_�	���޿�:T���,a�L┽:-Ҷ�HIK#u�hE��8>Ͻ�@_� ��GT}P@ �2{**��b��'����/����&#�a��6�ؓ�:��tP�ն���U_�x�6N?f%���hXz�bL�\ŷk��bǁ���T�˷��f��������ߛ5�����pt�$�_J;l'_��%E⓾l|w�x�&z}+�;4�s�\ƿ��=ƛ_myR��P����T��?ko9�~
�ǎ�b{S���FE�Ђ�f�JKK�W���`���}]g(��'����A&�{��י�i؀��d����:�1��:V�2��S�Db�d�	��v�[(yg��J
�t-���'���wD���Z2��|":��>�����Qg��6*d[�'�Hg��PS��O�^Ćap��� Y��b�^K�䷟d�Eք������VA��e��G}��O%%��4y����?$�g5��Veى����gi���t>Q�cTQU;�Hb�� ��-'㐤���|*$B�/��<��e���d$RL!E�I=���pe6�wR@ޑ��a�p���[��
}�$��o����5k��@���_��Q�p���0{�*�Q"aH-{-�T�K�=K�#�����%z^uj}��u�����ЖE,���3dqc/)�^�Q�7�;��߉���������.���N:��^�f�G BO;X����]��./�v�h��soP����'�;��lo�d��:��$	qh�y��L�	����?H�o�ۑ6��x��Rc��ǃ���G>=gq	-��{��A����ނ�[jē� �T�ӣ6�����q�J�FX��ף��fU:���?��w�sr$��]��d�B���J9R�?�x�k����`+�������ǌW��`�j�Q��a�Ɣ�Y���[��8J�O�� ކ]��ԢR���7E����~2+�������I�Nr��O~u���O��ێS��IQ�[�E!fs��<�㎊���H3){��&�����L���x��܉��>�	$}�����O�1D�ͨ�IU���zW��{�����2u��]O3��u.I.Þ��+�KPH^͸�q������8�Je�9e�d�����j�[��Z]�ͯzS^��g�F-:���U�X�a����Sfp����
=AYٔ	7COp��W�d,JJ���r�T��8����:�WFc\���sr��oz�MY;?��L���{��u�7��+��L�3�C��G�<����寒򵎣�� ���w�Y������w{�)�GK���R�D� 8_`�c��Q�o[��r)8��M@�3�������»���� t� 7���1�������fB���Q�����@x�0�߳��|.�,hL�`���ME�B�	P��{w���V�j�t�X�j�c6�[�?|��֍\�H9�Vs=�	�	���BM/���큖�;h?`81VaTZW��M����T��.�ݒD(��0�盰�N���X�>R�Ѱ��-�6U3�b�@�*R=e�<���~]���05��wFvw\k��2�5k��V�L$��~@7����j�]�y������Y��������"�66X�&���MV+�u�L�2��k�Q��"�6vv�����@(�e?Q	��񉐭��J���fS2$�eÝU����p�����q��k0���	ц]�����<1E��{n�	��Z��AP�s{� �L=�b���rW�<��~����>/�u�3о;9���3.�:^�d�$��+�9��!*��4�Iԫa#�k<����7��j0��R�:C����7�}�X�FF�$���f���.a0?�Z�W��
Y&��3/���jQ�KR��'�Mq�~1�}Y�`'�OX��Py`������2��/EC���W#������@VG�5y{�j��[<��}4yQ,+�_��L�;˦*���{(7e�hODc�R	���P"�O�!�|+`�7h��o�w�!=���.s�4vǄ�!ò��(��OL��2Ѯ{.a���R}���fy;2ݴ��e��[��l_��b ������D)/�e6�e��zT���آe%���q@Q���I�f�WQ��?ߵǔ���r���$%���9�k��V�d�w !߻�)@�����~���U����m���o���fgz��7��3��Z���"qta�RR��I###t�H����~U����'!)����������{�)>&�᝹:c�FN|2y�3p�z06	����"����B1̒y|��*�H�}���o�X�d���6��Ï˥��Wo�zuT{we���<����d��gJ:Q��'�/�"^�kf�N�v�c�+~���|*����^<l����v���.���m����dz1��Oѳ�'���]V�,�\���U��J��$�W3��5��3E��dOP���x�sV)�Ϥ$0;�yn�(C!�Yp�WN�t��=
*8|u�<픤o� �y�:��Ȩwa_�!^,�׉kp� ������ry�8��%�5�
���\:t�����R)Ļ�~�&�bT�L�V�"��_^h]d袞�Iv�S��B��Z_�2��#�>א01�mX�k���g�=+�<�p,��E;��@��w�����¸�/����I�O����k:�H�!�xZɀ��|�@�\SQ �lmm%db-�������|��\X ���f[�Fyr������#��V?�Lv�@o��������݆��a�{JL�tFz� ��Lg[�'����NN���M/��k��2�b�7t�h����,�E��S6��Z]����<klP�>v{�8`��=��O�E}rp�n�_�S��{�j����J�/B�iUu5؇��p$@�m-���I�)+v�=�X��Z�'�0O2s8���D�K���ۓ�m$�*�����F��O_z�O��\�Q��DI �* "�4H ��qɳy?^���]!C����py�uǽ���%߰^!QɄ��[[�)��ɓ�I�����Z����~5��4G�j3,��t�t�Y��O�F+������㟭k��cSS����a�p[q?��D3����+��Zfe�+�Z�fD�w6�s�`�a�[z<#�:�����
o��G�_�����G��#�Q�a�m�b'����%#�F�1�]*�)����A��'�!����0�����`۹)�����������7�!����]���*\h�U�)A�ɻ/e����l/�׫�����@<?#EUE�9�jaar�yy2�� --X�P�Z__���.�.��Kk����{�臾��x(|A��6�B���e��{���Ĥ���-!���G&��m/�_E���u��;�c`q�LM=�j��	�L����� K�/�n����S�s�ڔ����O��7�*$�j�!d��	�w���aL��'��,����C���O��c	5eN�R��D+��-�3%u��WM�\�8�F:�)z�zwjy1<����U)�U��9�o�����~a�{���y#��y�=�~�'����s��w��d�2V�9Lw���^Q $L-T����]���L�j�vޭ9)��^�P�Y;R^=
���:l���z������I��ex^75���~�Jb���������<0�E��O��{��꥚���ib\������;*�g,��\���ed +X����.�5�r�W������G�6��������/�R�G��~ɮ_�sx����0���d��r�@�6g���0b�h9����c`*�],��0�����3t]��#{w�'Gb����;��-k[eb#�4����\�A���gE�x��%�j��N\�������RM!f��&@��7�<�$pK��b��-�@xM�`V�0���r���崸�R�SO�1���y+o{��)K�����O�%�Nm�+E�3\dW�kΖ�i�=���=�n
��9d��R�i�jJ�r��Na�4��U���"4�#DN��9�#�krr=Fee�#�9NAA�Q��`Gb��L��ш4;<$d��#@�	���b	�}�����e���1�g2�)T�L��HRRk;'��r�Zh�0��<<2���9﫩����㽰;\ � pѦzu7��{m8����w�I0��_Ow6�=ǎ�/�l��F��F2M��p��^�ojf�^����mc�� 	���ڈ��F ��Xr����!��Px�/^�m�;�r�ca ^�� �<a�,���f�m��+ٴ��b�yMW>�xM{��N��HĐ$Y�O+��ɜ5��T���	�.~��S<t�%퍤���}����6_xmooW��3�AX�Ɔ��V�i>[y����v��7<|<Ai����7�4�h���Oϲp��jK��@��u���!;+�/f�/9������=��oE���>��ND!66�c�`pYX�-����.©�T��[@G\�d��S:F���}]����U�%2�5��W�:�`+�w/[ـ_�
'��G2�I�����͕�V�F�%b�Svo�agD$!a�0l����ޗ�L�z�$
��<\�{���!mԩ�F�93��|����T8�V{��C�]/��?۰�T���Q��B�LYYa��+�B�jy����T����M�G�	�#��֝��Zm��p�9�#�>G�wn��a,r�bs�X!#�=>�)�m@��c����%��B�����a� ���>�����)7��3���n�潕�k<�6���]+ߦ��O�Z��55�8�)Ē�l2��P��m7mG7��Z�Q�ЅfGRIIɲ��ψ�'E\D;�,b7��F���u��5fTy�^ASJ[
���]cϢą����5�9 �׭[�ݲE�g�)>dgZO��V�s=s~��_L�T�����w�K��R1=^DMB�1` ա��:SZ���S%%�|ji�z'�ak�U��}}F��el��;�"�D�/SI�~�-�������,���KD�j�}���
�ʕ��5�x���qy�O&�	k �v���g#��ԯvK�0O߻g���x��(Tl�U.O��W��c<{�����ASzG;Q�8�Jdo�}}�=���3��W����>��� T7���f�&`Q�/�]��"���8T�* {�E���Gc�f�z�CO/�>xv��/��8�{�ZUt�Ҍ&{:4:�ibb�>�TY����|Y���6*���-O�p�wm+;;��EC.�����45[UU�< ��yx��%��Dd�\��" l��E˙oqs3��R�M�K�E��pB��qo����s<tr6gz*���=�{����Nm.��W�L
#�Ap�D�1��&�H������㚏�1�gQ�p���Y���W����ܾ�Tl<C5�}�
�ׯ�(ʍ��C}�GU�|v���ztG�]f���i\O0�"���6�`�KLW�Qn�βC�綌sn��M!O,\�JDWk��R�S&��-�7��>hu�=�[�Y��&�ޯt�ȷ��ҺNgf���X1�s[J=[j5/̆� a�0���� ;�Y<X��8��ώ����T��B�;+T�[�`�-â�&6Z�"gqf�>������a�������Y�p��� R"ù+5c����c8�&A.�C8��Y�_��+�<�M�!�����@�p?�d)��.��v���������"N����j"�]�⌊���;;���I��|��ݩ������h���SWG����5`��Ğ:/|���	�;�k��#�3�(_@��B�@�u�����Lx��nq,y?��ο=(��6��iJ4�0�dp�.��Gk��\Ȇ����,ߣ���ӗ�o�L�n�Ok_�/[��4$ y�0�NǃZ�xR�������ӊ�f�.'!�{V������Kl������W�+�3��T�;/�魥X(�s7�yl����������ؖ�ص���,���n�w~2��U�����cXHt���
���Bd]uף� ���p�h�D�_B�V��m3[����OԎ�Q��������X��{�7�r�����i$����=Q������D�Ǜ�+D�f���;�lV�L�
m�D:xV'2�V�W���WC�����{�w���eb�/�������,y�0O��1h�Dʟy�(o��C��M���S����p�0��nQU�!pR�3f�8$?S �Y���_+�nIlf�o��B�"|5c(���_'o�aJ嶚8�N�9ԏ:@>2���(�鷰�8�z�����[m�7}�cr%=��k����Ӣk|II)F]�!d,���w�+�at�M�s�.2��5���VN` <t�pi��soមk[0����߫���ҧ�_�/1Z�����K
�X�����!�@~zs;Y�]Jŝ�#G��������i��C ��TTT����WR�'
���D����k+|&��L��f���M�ϵ�8�ͯ�04�Z�����l�m�x�M�l�/��^fe������;�e�\ާ�;}���z���i��zB���?�O��z O��Wi!�i�}V�c�8V]九-�1�_'i�Lj}CA��!�;� �}]%ů�\�Y�=3��9��n�j����Q]�*�����G�}�F9C��q }���T.AF�'ȃyڃ�p�_�F'���O׮���Y�r-�vҠ|�3z��&,%������J[3�IVN�8��b�ޱHh}��n��dG�u�7�+}h'`&��հ���SA��c�R#������Z�@\�&�g��F�c�[;lv�Uƾ�_ 4(�B�oY&����F�:��ޖ6�ܖ7E�܇:�M=9�ȏ���`�GL���T�9tI)��M.����w&���F���nM�u����x���gAPWbA�e�3_�d[�t\��O�c0�y��ɬ��T���g�j�M���Z�P�������Y������X�`kW����Ŵ=��v�^�9�z���u�l�R�^ژ�����%�U҈��d�#�q���n,��oP��G��ƍ�����j���Eg�n�<aŕ� y����c� `���v,���2����&���{.K�E��q��'F���2��8L> �p'*8LqN���1�*5g_Î���<��}[���
����,��=x��1P�&eb���[y������`{H���ac#L7����'��饈>����.�XTi���Sצg96yz�ƓP���[Խ�>o֯{�`pi_�#
��j�����\ScRXt��6�s�=���$۾�f�8j��SƸľe3�F��Η�S�Ь���"q%�?�@yE��b�B5 4O���IBϥ�Y��刯`����{���U���� �F���t���/l�J�قf�^��s��2�L]��H����/o�t��|-���(L������дq�^��4�U�?J�gy*�μ�}`�W�|5zKmcbc�Ng�ĩ��) {���p�r�i^��:�=��9� ��IJ�ZQ=lԩ�<��>�pʯ1'�b���x1TSF�O�3��)��}�kОM�����R�?��'/t�r��7Ęo���S\�ש ��E{�ԯ~
{�����w�@���G�2��N8X�:X�"���'6vKO~���U�۝�d�^�����)�.�d4�o��/��ܖ��'�^0bE��e�[��fl�!H���7�ӏ�[���z:n5��7M��H�r�vk��;�����{��� 'Veoo�����a�_O%&|�9- ({�;��^�v<*��{�Z�
S=����ݓ)���n,������Y�ۻO|"���AE�WB!ɇ�h��#��w���c�ںl_Ӻ�m�R׶��@?�ig��%G�X��U�pG����ZK���#+?~Q��S.� ���AS q9.dH�����H���ݛ�o���|���@p�,I�{)O�?DN���8�I�ox_8�0�=w7G�eevoM���wM�x7>�W�<�=�Y�������b��'�grl�,2(�3��::����c"��:<�yF�C���o�0]�!ߟ�\��	=���!6G�/�rFq��Oh�Z���a��TG��g9sT���[��9��Ɍ��*�rm�tC&��z�[���a`����	�q�Q�P��)���|�k��{�p�6�tg�z�����+�`>pw}�
�z��gNO�z-A����>��HtTvR-�n�� �j���Ĥ���:���m�ٖH�~��8(���'Se
R��Fz�e(-ZR[$�YP��`T�I%�u3P>Uu�2,��xb�_P$��\���U�A�N}����&�/�>�a�Y	:*��Yy����kۛG���(�¼������۷��JY]�l�9��h�|f��&��Y6�2�wq�8���ĚK�"\&���ߩ�^�������=*�u��N�E]�E�@�����ͽ%>'�FVo|�U�{��o/m<ݲ�_�Ϩl@|�2#��yĊ�v�N��!���:���O�Nt�4���Z�\����wkFB�Н���=�;�t�C���E�C�����������:mtz�Ɖ{���mh'���C�\7��Aq��wؐ�������;5���y�\D�?G�kQ!�޻Ab�6���j, t4U5	�(h���_���	�pHߺ�1����	��Խj�b8r����+z2�GEA�p�H����s�Xs]��}�gR�mPG��m��s�n�B�������ϟ�m���9�op��$.�y����ָ坠L4�Fx�e9X�F�hq�ӈ��vɴL7%�v�/Ci�� �~>�-:t�^d�Q�HS��[ʑݧ������_��B�8��i����Ȍp�黿��^`���N�4�VR��U�#ď���8<�)+�vIe�O}=�q��8,���A��#�#��V`וM�xH+#����A�R��z����y��L�Ċ��]4x�9��ږ���uG�E�ތVg�7��8���$ r�螯?{'��6�|;[�cP.��(��h��/�j�oku��
d�T�}����m�����3���I/M�{Tz��)�?� ��3�Q�-�Ɵ�A2���i�
� z��)����PMOg��&I�a[/��_��g�|[,������p�.6!�Ch���x ���D�`����B��cߧ��'s!O�{[kʩ�:ɞ�=/	\���vJ�����M��}b����z���ug@?�NB�ރi!�ߖ�U���<g���v:���/�m�݌I&�u��充[|��0)�4��(�~LП%Ŏ5��F&?DxG
Lo������].{p���V���WٟxcX�j�ƝTQ��b� �П�X3%�V �3�8�&<Zk�D�,���l�uT�{rd�DY�� {V������2���|N]�k8�u�(*��[#�����zqj�&��a2�y����isr��W���Ϗ)P�1e�U�����g/w�?����LR��(���2d�����C��_2�Q��T0J	w�h¼������~�x�v=24�r��EC{�����w.��{�P��������+�$���Y���ӎgY�:>��ue��¶1՛1�"�^���%\~Ad"�7]#�ȭ(���	1��~ݴ;�
�ZI����5��]E� ��]'6_X�AY�=�|U0��d��:���݀��i5O2��O���[NE�ZY*8׎��/�:��a�
����WЀ������[�z�O�SLI�w�}B����c44vx닐r2/�Z	5�*�^R)~����~�����R�=�G)q���o����{���=*$��_5i"�7�-%goܗ����lr�KN�����Z ȗ����t6M&���) Dǰ�U8ER�-�`�ߠ��񫷟o�m�g�Q�2ӳ���8C@�AA�@
z��H(s�Q�W0Ц��	He�� ű��BU$�Z֚��U@���_<���p{�(���N�ޅ�CKwO3�G*�1W5���A�&E�������)�������kL>�D�,5&��z�{�-6�^�>YC2�w���,�×[eP�mfoǢ�
1Bd��:��?���~L�OKVnؤ�U�E]���܃m+s�0��L�<�����3&�7�i������Ͼ�x^����j�&k]���|��>$h�+y~мS�qp*����T�@�m0:JЇ��2���[��)�kM~���B���yG�M���M#�����B���(٭-�ɋb�e-U?�{%���V��\�.=;��m�����2~�T��~<��L$�g\8���Z^�69L�M��c�B�I�]#��!m#�σ��)3_����vE�lk����q8س��jV{�\ʱ2��+��x�.��������K{�Iar�ĝA��B��1���l�_H�+�ф�곲^=1b�`�c��_������6� ��/X>�V��Uv��-o�x"4����4���&)3n��(d��B�z5�>s�za-�n���&gq?<�yI ���ɳ�#W�H}v��p�V��i�W�_}���99��n������tϭ�I�{�~��t%+{P�u�V/M�t��4��w�������S�ᢹ��b�4,�S��^����n7�鵫�R!��?��M�|���Jm�Rf06���{C�s�4iD��=d�6�|�sص�T|f�Yh�ޒf��K�+ف��|�{�O5ܡ"�?uv.�߼>h7��p�Jr8�Q���<��$����i�7���_��J�E�ռ��c<�	Y��V�H?6��5� 4|�$s��X� U��#W
�)c_t��8I"vū� ��G�XM�쇮Qoh��\k	���;��Q�.���@��.d�2�߯l3���e�����UkM3*F˸����`��wΥ]@����G��;����o�Lw�������v�k�I!�1���;ˊ\�hS��j��<,�R�p�N�e��Ƈ��˖R�0��!��}��Q$��[���Z�y��ҭ�8�r}����0��mʤ�@y�Q�/Q� ���q��c;�)�9>b�gP����މq��
C�l~��d���d�i�6��W�=����m��c���Ο>|f��ܬ����_���7��kDav�)ᵅ���g��BBdzN���h�ke#�7����m�\c����F)��g��WU�(�'��:��+;@4��QK>�[^�d�Ur'�l,�N���mp9iߗ�c!�^lc���E:��D0u��@<eS!j�o�0L� h̀c��_91���	w\��  ��Y�H��z='�ZH��n��|Oh�`nr�yr��^�nHҐ����W��*^A`O�l�Ƕ,�pCyEMQ ���~��5�կ~�Q\��[� <!^��a�y��|y��)�b.�.-��"?���%�e���z��� 5���V;{~*8���
FBW[��S=@�3J'���U�	��}��YZ����0w��l$t�y�q�b�>�B�@��X��+�m��}]T��M)X��K���r���h��|���Q���{��g<�ʝ
�k��A�>7��)QN�V&�ט��>�N���C%%�)sn��wk+|чK|�jٔ��f.�J[�ЎUe0��a�������>n�q"���pws�Py;vwE;<2�-��ϟ�^_�ȩv�F���e�O,�~�������#�ͲX(4*����k�"�@���������f7Ə�K %�G��jumF�/���3��/;s�Hŝ:N����|,�/��E�s���~�?�����ō���L�4l4���L�Vq��t%��P�q��W:`�x[q��.�&~dY��yՔϚ/IL��5��T�x �"}��/^�����.y�%�fZ�s\�Hp %�	�>,��Z�yk���ׅ��2�4ǡ�|�?"({>  +a�=q��H������P��zJCf"�nj[�5;�;?�J(�m��ƫS������?1�#�
�#����`��+��G~��5|!2����x�r��Tɱ��tƍ
\8���lw��R�͢���є���m��DVN
G�;�kg��q�	�s��\/E'�(�q�RΦ=��7Mr~]+G���?J[T%�7n��{��$�3e͐>�k�q����7��b�2����iW�]�(�⠳\�m" ɗ����߹�7Z���F� �+j�(l��c��j��L0Nxt�4�`��o4q�ڦ>�¬�q)l@D@�FqM�zA֚���(�\��eG:�{վ��30��Tx�{_p���wE���X�*(q�kW󽅳cU�r���ٿ�
Mʞ��*��	NF��`������F������dd���n����eP����w�S��߁@GQ��:UW�����������)	�Z���x5%bfG4�5A�!8CeN�~��?�z���υ궊2P��;F՛�7��vN�����<�����L��I[^q��tKATv{���'[�iF�i�,YF���`Sח�ɏv&���rOt�X?��aLa�t]*d�l0Zv�W��A�A�L�L�`��:ڤ(P��~nE�v��1;�&6���J��r"
�`n�T.�u�}�k&Ch>�*�k��e�U;+EqS�Ǐ".B��2?d !BN?�;V����2y���W���U��>���q6�qy�1���<�\�0�n�aLaWgv�q����9�����.}]!����\}r��)ͣ���=��j����R��	�V(=f<�k�fA�n��Ι.�U�D]^C$)$��o��{_MlL�dwJ8h���F�jia�mu�j���Z�2��>����F��^`�9rPӇ]����*�
�1]B�a�������Lj��f�:AI��ON$��6}m�&d��
�u�*s������cb� Qo�t�����R��$�f(��Aa���o�j�+M5�*�oh�U�g6��jk��qZM�?�f�O���M�������'�F�s�Y7͵�8�_����jܶ�V�G���ݡQ@����������h�6���>���6�={�u}2�2�K�U&�����bE��F2�%�.�-W�I�Y��dDK[�֭��1u��r�u��Q��և�||:c��/py䵚�ij��=���+�A���]'	��2��#�krX������e�_���-����u�,!m���(���(�����!R�aYki�kly�'ü}bT�������c��7u�'��D��	�ix%��+�Sk��&� )�f�&�*(&%�F?k^�HD&�Y3B�qtys �e1���|n����®�����o�1��+��;ٗjj�{X�c�⟏0\���)^�T�̗/� ����rW����Q�D�$�n����}���m����D֋��O���k������X6�����(g���<�����l�]?���4��O�X�k˶
��0����E��q������?Ǫ��C^L�엔����FU-H���y��thp�?9�W���.��B�>o�qb��������j@�f�p�]A�� DC�����`���x���ync�z6������y�4��_.ڔ���{6��a�8"Q�L��#��/#��Q�I`
��g/��������<q�I������������^�a7~f/�g<�Pƽh�=��-������T/&����u��z}�C��J��'��?�+���#��o�JT>e������m�R�r�[�}U]MU�i7���U떕d�&S�����C|���~�T�]Џ�?	���)�r�7�4x1��������~QD�yB��i3+�fd)��C�;�	�݀E��,i` �s���{i��7��?[je$<S���cY�`U�׿��*׿��c��9��*{�aV�.!0J�g#�L�V��c:�G�**\��(^o��(�հ�US�J��I� uoE>�	�F� ��f����ui�h���o�q"ZחE�h��ZK�΢+��&�������T�-⫔�1k�K��S������>��78�lvll��'�ITܔ�u���}���TK�fvl�HE@Q5��d	5
o�d����5�kQ�֔�Rq&`)��mT������ݗ��u��w�{��J�q�7R��A����X�7%�� Zz�������2��8o�ɻ�]C}j Ǌߋa�hqF%$$Ե�+<
����i_�wIGU�\�!^ғ�M�
{�~0��uB��඗+����T��a����$L/g�3�a��X��� FھokZ�N�n�K�A���$J�v\�n�l�� ��KGf����{��2=�S6t4���u��Ń6>܈2��t���~�<IBdtt��،ŏ%;$|����a��'#{k�@JW�C���غ��?  � �a�Aʹ�R�1YEPX �����K�6|��A�f�\�G��J�����:<�.@��-^KpY�%oou�]ng�&�����w'v�ݿ�'�U�ї�CA��?�[�/%��.�f��^amc߯�oŋ�ABT����15%_>2	�3��`�h\x������/��;^͓������ZJ=#��\��8NK��`oio�h�F��y�+�8Ō2{��"5Z_�(%������}�d�;H �ʞQj�M�;�4���n�Q_����a7��~��|�3��Ia���\���ݻ��Y~�^��✻��W�UWa�ə#�\�ee {zz�V�n�>����G�)����i6P��	@���T~m�BP���ؾ�u���2+`#n Aw{��;���ш_�$2�W��+��X��!毷V/��uK�*q��jެ��費-���.5Yc�0JF��-{1B�
��=|EIIY�o������@�:Y�U�<�Ƣ�m0�2����CL�Cp�mlR����>௦!<�����y�=+Ǵ�QE���zd�� c���:�=��9_�������G*�H}���q��������L]��͹���l�|���z�k��~\���¯�uݒ>׏�;��S������M��ׅۢj�ޔZ5kojU�Q#j����U�gѢZ��,�v��{� �.�D����}�?�~����9��s�9J=_
��q^q!Gf���*Z�_~��W)�CѺ_�-�&$$+�ᨊ�<��i.��8Ǵ�����xs����E{���G�Ը�{,�Խ6y�T�D�W7d圣KA�/���[Q�@��P!��b�Dv�|��~Eyu5"����ۯP��ײ��~����K���Ŵ����觸$6��½(�5��pu-Wп;0<� ap����ϧ��e�Lbu�v���ͺ���e���v���X�#pBh�zlNWق,����O�|�G8
�G�9����Rc7����X�4���uz��Qg��8L�:��*��N����p��PG껕�3Û?ĎX�i��f�"K?���m�J��cLzx}�t��G���2�q��L�-��7�_�PG�����x���0�~-,Th������\���SSs�{'`w����b��aT��b>J*����0g̕�>�es�zaR��#�t'a3�j��N$i���T�mG��>�l�yZ.�� $��z�*�����s�2A�#˕){�X��9]��͘��d�[OHO������AU\�ԁ�I�e�v�<$����2?�����9G�A���R�:��+-$�^�X��������7t��N�v�./���!gڰG_>��>RF\�}�.Q�u��Ӣ�><�&�����a4��f�����KV�l}�TCBҶ"�la�.(�nڤ��%+�n,�~{
[�=^7a)D��L���%?���;}�s���yHQ{E�D"7.��lc�T劌����=4�E4����ަ��>m�F $�n-P� ��c��!�b���r�������)�g��d��~�������踮gl�Z�"h�iQ'R�Iԭ�Z�
H
�g�	��ҥ������7���_�/E��͊��\Fl1%�O�Uf���gS6I��[CZ��}je9.�S�����J-�P��ƛ.�(:L;��E��J:����*�X��^��x�5���Zb�e`U2�l)���T�봸����c����O���/`�:�z�I��������c=B橨����(����g�Wxڟ�$�/H�gK���ݘ�Urjm�L���#gu
��m_��[?��|��[!hZ=NNi1zq��|X72����"y�*���K|��@\�t��?T1��	�s0ӝ���3��'f/2�}g�ZI��K�2�/C�V�"r���d���#l�d����P홍��Y��lgL	���ψI1t^��z]�^zeQ��,!�j����(�k�a�,V|��˨����Q]
� �N��C���*����S�D�����	���s�Z��}��ɟD)jG������S�&�}qs����y��3�
�.���'�A4h����`�j[�k����±`�E��M$�d.�R�����x��B랉S��Fe|+z�����lڂ:E�`�X �qa��g�&�/;���~"/Y����P��{�w�8��fk��yB^N�z����������u��Ie����^���D�����?��66��L�sb꭭n�c�ЪZ�oEd#8+��oڭ��;(��&H̀�;��O�T��
`Ig�2�#J����H��Z� ܰ��:��%������[��z��L|�#��ϫ�N���%D��{�y��jIF����1����oEzb#�l��:�6q���>\�_��`���ߋLD���nC��uk��0�O��.J|�U)J;#n��:��8Զs
���r'ӑ'�/{To�iڐ|���������!���xGT�秠��)~o�DV[���}W��߈�k���1�����sttD1���E^��3��X��y��X�=Lc{�K	��Cvs����#�輻�3;���j2�>k�����`|h���Y2s����KT��+��ȂuJ�4-�[��$Ҍ\j�r��O]�]d�w���!�XVyZlEf���'\��L=��;�q���.cOg���������Oš���.�-��̜-`�"�b�8b�C���q���C�4�B���8;Z���;��f�烼WG)�+�ߋ��L�o�� �<h�{�Iԅ
����cS'w°t�:�N�tu�@j����xsj^<R����D?��� ���W��Y�c����o�'u��
b:ְ���C����۫ߥ�)̷Ǳ)���ψ<�޼���WYƔG��C|��:/�|���U1��[�������8G�z�����o���F���C �J܍�]�
r����F�����k�>��
���'�*��-�J���\&���<��OM?,�38u�e��]E�z�o<j���q�<cˤ��<{Y�]��y���������
l�<���#z�̼b�.�*�x�p�����,�|rK:���:r��]2�+ɓ���K�|@@������S��X���co��j�9�.s��r�)�-�ފ�12������6�a�>������ǫ�v����^֓���K5KtV�������}�pY��?��	���_��y �w�ܤ��.4��{�Zyؔ��ύ0�+��	�<���jĥ42�X����8e�$��ڕ�n�?�l�-%[���֗��I���g.aN�C�_Z��J�Ը;�b1�x<�O�j�e������(�]~ki���WQRz��[�)`��q$S)k)d��|���!gD�0o<]�dwߒ����f���&иf�ēBpڂ�{d���o��U������"���=@�}	��T���=
�s�a0.�)���Ϭ�E(�CNc	�2�ٵ�}���?���:t�DəC����nm�K�<F���0�Y�$ä4��#W?	;H��T$&Yi�_`���'<k/ŗo
"�_0�x��@��<`Y�e/�7G�B��;�/�̷#F���j.Y2h�������6�W͏���ql�k�3�"ޚ��*�)n=�hf�����mI�}ڷ�I ��~���t��������O���������b>N6�֮Yhz�9��vY��9�"�6���7S�'���b�K��C��Ta��魍��=�q����J��h��A�?�5��X�z�,�BH/�^�qD���q�c������C�^�U��Wm���|]�4PGl �hF8����n耒}�i�Lo���G�=4�6ؘ��I��lnT��oG�d��4�oE|LA��Ӵ���.�i��2��(M���ֺGQ4��Ҡ(�eyRo~5a�?˿���0^��\n�+HJwW��_R�Z9`"2ob/���$y
9,�,2~��OnO�m�X��PY����7��Xg�RR7-�n5|���-��_hp�"Y.������L��IQ	()�?s$
M+iL.�_]@���Z�֬Q��u�>%.��4-]���&:(��T�6��T��xY='�S���OP���{�7�ǥ��vV����j8���97t/�hyς*��8��5�m�h�����E4��d���c��h�ѹV|*����G
�w!�$�͗�Õ�{���YX�Vp��&�
�pe-�PDs0p������O6cIp D�R.�(dN��i� ����J�����*S�����!-��䬸1�x�f$��@�mP�<j����%`%(e3}so���������d��<^[�S�N�q�(�:�`N�E�� /�T���/Q#�Fd��G��vա�_K!��T}i�bџ���������ة�y'�
�~r����d5�%��e��F|z^&u����Y����@�ި������YKk�i�6?͙q�x�]�/^S�`��0[
L�/�����* SS�¡�����%^՛6�\F����͗�1�CÂ�(ɦ������%���O�\0�v�A�R�����ӿtc�S1U��P�o���&�r��(PF��*>i�շ��!ۘO���+
�9��ח����
:$�mM�̡���_&��-$`R�f��k]7j_�\�5Ñ1�g������R��[	�gۥ�q	V��ϡYq�!H�9؟P%��2y�Y���~ȺY��OW�vX�xBG��|-T�tY�;���G�l�q��O$�թ��l���Ӝ�l��C{���'�ԢeK�9���f�
x��OAa��Ѝ���)�/X ���4�?H�eJ�r��������� b�#�9��A�[mW>w+1E��u��;��g^�
�q�\��{9����������|���M�' ƛ̈́�u��񞰣Q�^Y���c�b)�Dě�p��E�9ju�GsE�=�B�S~��Wى\�l������m�Հ�HG�In��,!k�f�b�#�v�cӒ}�� m��ju {Vw]z�/qu�NN��&����ZE��O�?���� v��-�k�mC|Y����[�G儙�e
m�f�+��� ��X�N�$������I^A�ӊ76JJX���'�������~�`��G|+�DC�8n��8����Ֆܦ�,N��秒��M�Mw�(�������=�3��-��g{���{��ʞ��bhʤFj�y����r4��obAhf���/��ux]��(�����<Js�]}�2�WQ2r���`#�a�HK���-�^�Z\dpԽS��k�?1�
2ϫ���lu���a���v	6#�C�{���3w֚�Tª�}�j��4�.E5�u��y^� ~FjlĎh�L��n�ΞI" ��,�^�ǥ�]n��d-6�F�~�$����xX�=�^e�dI![4k�3�&(#���πIv�8�Q��:�)->��T�-�Z�h�d{ZFq��T�M����J���je--"��Kk�OB%l����u�N��`�s�$��YKy���Jz��j�R�S�WU���TQ�)��9�S�ߊ��H�3�����f�P��IS~����"	��h��@�o�|�u�_کljj�h)`=�Y�w�}���^��|
 	�^�|G�ȍ}�݌��m�z��]>�D$�����\�СN�ͪ����'_�q�?y�vE䓁DV�6���K��vYHk�ݗl�"'��+	���hgE<%H�F��p�a��}/���ɷY��7��-���������V�����e�����w�{����������M/��?z���j�{;���¯K���&ce����[����s���)�+T��G5�� ռ/<�8���u�T�a�U���g��5=�zWQ��s��Z�9�XH���΃�z�\	�=�\q#��it�^��=a�H��_H�j�1���n�s��(�2��O���B��i3���iT$n��G��л�hʟ8Dl�l�sq/���.���t�U!}ι/.�M�|���2��L�R1���6$b]��vN��Aǅ��S|�4�� ���
�� �=���H���v���[���b̕���1����~^Q���N> p��F6!�x���җ�:�L�r��ԟGȽ�ԩ�R3�� �`��8 �0�nz��;��6@�Z)��NR�m;QNf��~,�ޖ��ھ�dY_x��B���sDD=��W�5�t��D`�u=��I���;_�E	�,���ܚHk�8���ӗ�/�4Z�ih���齌'G�.��PH-.���M~���]hl*z�_s�]kR����O�ݞ�>�L�#�I�k&�-+#b
�}�����Cٔp�5eZ?k����5�׆{��[C{���i-�ʶ���as׷���V����kYJBε(��g�J�DFPo  G/=<jꙋ[��=a�.!���H���;E+��=�WKL��٣����Bo���Vu"��nq)�4t,)L�#Q]W(��ks�8��Ӹ���z���i�2��&�4 �e�E"@�ϝ^T��y�#7���D�<;���ˮ�Q�`;���K�`3l�^��<��̉Y^�s�w���A��k��%_�=�a +��o��%<��Wh/���LE�����
>�o�xE{4�t'h��1/��Z����R!���LY�
<��_4&����2{O�y���x���+��Wl���G[�d����kA����$�]UX�+�%���^��H&��D_��E�Ć9��2�E��qHcu�]��xT�"hY�i���s�ՀvL�It����f`jʟ�r��5|�uN.[�����.!0���Gy�ܡ+вE���A�����;,�!�^�7e�b
yI0em�]5����qU���E/��Iy�R�t|�{̣A��pW8Q~tt� 3�{+!�T�0Ǚ-ݯ	W^�G���<�0\A1_���/��1��})��eNqFb��9���jo��
���p���#:oKO-}���>��76�-8G��͹� ������w�$�
by��L�]݆��g<M����A��o�4E�)S�q�&2bx9	�y����w���0&0�3`X�r�u���H�V L������U�֔�9��)$�6��qSKKIL ¯���C�ʵꯛ������� �@^Ycy^��9��F���Nq}@�_�ܹ,�	ڽ�x�����K}�r��;���qdFF�Ѽ�����( �*�aYZ�$�|�G���%��j����#��'�(�<�O������yq���N*�%hմ�[`�n�番���|�y����G��¡�ЕX�omr��������OH�=WH��v�d������aA��aQ<l�Op�N^zn����n<1����2�?.���|�!�C��N�gi.�m�XF2O�
���+��Z�xA/H��s��҇������v��Q�^��=�5���r�g;c�*���o�	���X����~+���P���C0�-x�@"�籶�͟WD�	^hu0�^w�kV�M*!0c@k� Z���������S�(�q9>�UͿg�Q��O�M��(��cm���.�wy������F5?��`���|�f� �,<�� 6՚:�=�'�2hn��'B��[9�$tRy�NW!��t���8�:�|B����` �^,Qߐ�;����ѣ�F����3��]��ʡ��C��D��c䈙�[�톿u��xA�#ALK�;��Ñu:�à\�Q�N�����j��U�P�g��a��;crON�d��K,+^�,���p�b����.n�z
f��I��E�y����a�U;8!�N�H�o9�����X��ёF�w1��Å^c�Pe�Cg��G���R�^�����n`�L{��!3Z��P����K��lT?HU��^Z-�Z�E(���wg�Y��@Ҝf+�����A���0OBQ�
`RI��2G�����n<��R��G[Ӵ��6��>�c���
3���R)�%�
��C��J݇�R�3����'o\S����0�-?:fw{�q�ס6s�ς[A�,~�K�����NN�!鎓7�L=p�4�"Z�j�A&�˟A�/���fW1�4�v�O��]�d�<���ݧ���xm:���9��^o~�X����*l����,K��v�z�`4������H�j_��`��\����#���m��Z����r����@�,[�PD�S������G�O�/�.+�䀤{��@�j�^�iW�N��n�MY�UN�Eƣ��'����|�m;9�A�c���q��d�ۆ������^mx�V���4b��'��O/��O<�������x��<�n>�]t�L���<�Z��G��-��j���S��_m�x����W�^��E�t<�'���ł4Bz�z�-Ɗ���~Pы��}�P�!1sO��-h����վ�WA����wz�xk9ˋ5����-��
��=���2#�r:�H� ��C�SȎΘ]w��c�$�T�����-����2b�#�O�_I�d�Ҡ,�O0Ζ��;/סLb�ō~���~Do7��x�R�ٸ4	�ͩ�0	И�!k/xD�Rb{��Ίm 3U�E>۶H5�Gm~����9@i��G���� u�͋�� �����侂
�_ BA��ohƜ��.�9P�v���B���a!���h��E4-w<	6�����F�V/�r:�?{x�Z>�a�t4��Bs�c�%e�*ww}����y�*>�C���YsJ��?�\9�5��"���ʺ���姀�]���7T��w���?�s��`2���U���V7Hhf��<�VΘ�:�����!�n:��^��n�Np��9c.���Ϸ1 �2�X0�7�7�Ь�XJ�}�Q�Y5�χ��[�T�jܥ����U����_�ks��k�?C��pDGWF�5�T�*���[�!eF�0T��{����� L�����ހHDkd��u�s���s�o�PbQ%C�2�}��O�����/��,.XHc�+��������_�p�z����70rR>�W��I��p��p�/�C�3ه�)2Qv�f~�9�ɭ��#���83�2�
��3~��D/N�*s��e
�����a�/h��@T���mg���wڄ%X߹������(@��L��`�5B�z�%	���KG�E�|�$q[F,vZFCdF&H����l߅ �;7=�l�\/T ��PЎQ	�{m��@JV�w��"G�p�ۮ��]Z��j|�W��ъ'��m (��]�G;H��2����D$hj�>����Eܗ=����+�/L<f�ct��T�D�GlW�ѕA����ס���Ն��!��E�&_lKF�u|G��8j�|˖X�Zt��&yGE�Q�G���yB�n���l�@�nބ��O�[v�hP+�E��)�I�D���a�g譂G�=S�xE�}�&�H3��J%�O��*���]��\k�Y�o��6np&͟@�\?*L�&�)8���E�RG����a�2X�>/(��2:�	)��|G>o3;	z���8�KlvF?�A�T�k���/���jI܏�]���x��p�׼Z3����U��<�M|#�~�mV�.��	{`�쮊�iӇh!K9�����y�X���%�Ϛ��+�1g�5!%2�,S��s�Kd�_c_��>OHK�:6����`v����|�h�F�e}�����}�횙88�"q����zw���Gd����g��	!�p�"��w��"��@k�(��p�m�=::�=j�'"�^�M<M��\\�����&i�"v�K�̌g�`x6��l���*+2+ƾ�͘ʵ����l���^W[݈/#+z^��dN*�/�1.�M����?(����l��DD�i9��I��j~r��.D���!n�#�N>�����P�o�nTC�n��1�k���WPU�OI�z��x�F����U/�c��/��	<ÍT��ւN`��{���2�=_�������^���<(G缈s\.wN�zw����L/5�i��5:����V/dΙ(�ƈXo?�1q�o�=;�����6��=���j��������r[',���-�c��'w��9��_05
m4�'�D�է��6��6v�U:�!���K��Пջ
*[��q,�3��0��*D�q~����V�QU`� ��\z5sD�0i���t�ș��������M��uj<d�Z�d���]rL>>�:j���0��(V�/,��ܥJ�yc#BM*�MA�#'��+�;0�6���[��l$`u1Jdz��2���d'��T����3��~�3�9Ӻ�޲M{��;y������:�C��%����6y0US�H}P��9S����m�����������L��c�贛���n�r��~�j���u7d_(�Τuq8R�c�[J7�#����+0���S�K�ĒtG��@7��K;k��Θ�Kjxc2�sQ�^=^3��q �4���e�-�>����/{�<��H��<�؊��q<Czg�H��9�2?��m�E#�R)�V=qN����T�4#���|�m�M���2�׳f��u�Xr�ַ�F��Q�Ƥٺ%�?^N���[�鄓�^��"�w��^���{R��P�mi?b���"f��+W,TR�M�-Iyko��#8�q�ܓ�{X,�g2�cE�O��ԥ�����hl�,$���*8l�[����~�B+��h�����ᖖh�#�Ass��Åjd9Z���\�VyTN����Ok$�ǎ�?��hd@��6�c%��%�K��cKS4g��M���_��x�AM�������y%%U
o��~yw����'בy���p�jF�����-b����毗=1��%ԟ��4�k����sJg�X��i������ͷ��@\���e�����Eh{(��/�X�9%�#a�a��i5Aɗ{.�M[���U����4���gB�O>[	�t���\�
�4��r ԑb}ހd��o�2����g�Ś�u1��ؗ��$B̜WI��.��
�u�2�<��E�tw�������XonX���Pe��a?vB��k��2����\��ꡃѪ]���<-�6]�8e߿�-ʺ	6&N�[��q
ۃS�b 鋅~K��bޢ�=�> �ݵ�Z���~JD�KjjAG��{��6�|�d�i�*p{���g��
h�E�_�a頬�/�2�(vl��������߾��X�:�W�r���ү�^k)���H(��bu��k��5je�Z�\e�zsX�,e�O�nѣz�}dݼ����4�1|��t�ǩ��~B�&u|���/��_��J��,��~W�6�՘�M	*TP�W��Hw~��%T�FDw�#gt�� =F�כ*�>��2�l�_o�F� ���~��ʏX���w�I�����SA�
���u\�����}��hB���˶�sh/�	������kF,CpT���9���xB��� e��X-��r3�go*z�nN�Kq�)�ѧ�}� �?Oܳ�Nu�`d����u��J?��!�eaz=VnPQ0(������i7?@�!���%noJ�܌��e�yk(:��`\���9�d���r��-�����i�.eޘ���	THS��qx�kX�����2�im$�LƦLý!��ݙ
hm4�G�r�X�>��TJ�k�.�l^���D������Q�2W����nN1�wj��ё�]�>2-^1|�l��W���$Z��6RP�8戮��Y�
��2���Zǉ_�I��8�b�s�|�yj�~.�	<wH�SڱϞxd_�9we�A�9@�9�$찑�ʤ ~uA�:��V�����.[��Ꞔ������Q�4u���gXt��`�uE�|�v�sy�>��l��NNaBT9훾Xf]j�h���dߛ�J�%W�LoYq�QL��6����M��V��7��O/܇�R�9�6�B��#�)`ErL~B�ґ^8rێ:�̿e�5���Gͤ��u�h�*.�6
y�V_t�P�TG��Y73w�����hM5���2|H��$�Q��W 56���t��ڀ�jȔ�,RY�J_q�����1�즿�����l�ighZ��H139�`�����ԈVQ'SYq�h��5Nn����k���e��Aj��ҳ���)�����p���[Z_��p:��Sų�a?�w�@!xѯ�~x@�xA'vw[��f}�Z�W��6�2��=��5*����TIpn/��_8I���ZI��LiPJ[y-�����x��|W��\���\�H|�KD�9��yc�+g�t�� J��Zv�V؆qW��y����-�{N��5���B����N�{Y����a��>��=�����l�^�R�� WS�����Z��a'�"Y�U�����Un"G����5V(\��0*"��{h���[�^�ֳ`ꜫ��'S�/PCy)<W�9�O��
��p���!z �8<�A.�q%>�D	2U�H�{_/ �������1��uU|7�H���W������][CD��������_X�~ӽ(���VL���hڹo;��t��%bs��ْɚ/��{�8��?�y�׷��2=�`��r����, ���M�'R姹�;����O*�2�K�5�����T����bSM����o#��[5����3qɌΉ��j�-�-�9��ֹ9P�Ef�BMҧ5�����hfJ�?&�p��ï0j@_�&�=�˺z�\	�U�����i�b���)=͍��<�a����ӆ�&fyw��<�������:�j[�8��%
�W�aJi�}�]W"S�/�#I{�1�w
���H��i�#X�36(Q��5�g��;��MS��S�.��[�i��^�17>�*�W�q�pz��'���2����O�J��򴴟��9���߯��W��1Rp�_~�e��Y�/����b�/UUq�<V[r��~�J�]|�A�7�����r��s��x��w W2v�N�OZ�������"H�#c��9^����'ph{��`�u�2pk��s����v��*[L�|h����C?��S�.��
���Jf�L����L�w����1��_�\e�t���Y�XU&�pkA�O��;))8��)(i�LBg>ǟ��*v(CE�Ӈ�P%��i�F��⁁�v0Bvyy��� V(/"@���v6����q��;"3�J椗�F>,�M�SغQ�c��3�dӈ��a��9��x�}!�0�镣��C�"9%/L�n@�+�!Z�s�È�Ǿĭ4n�}R�c���Q��ĥ���ޗp�R���Αډ��J����X�P�N
��B������m��<�>��:ZZDttt2}ԟ��nz�2��Ne�|��'Wn$�%�勑%'ߋȫvg��,c�'�!�n:�,^���X����r�)�I(,q����b꩏ÞT���������[_)"�":ucߣP��E����B�دǐ�6G��ˇ��N-�l�*�I�E8;;OJ�S��8����������y�?�����)�Y02�P�]�
�����u���1B^��m��}��k�NWz.E�:j�~m��@^>+s[uS�oii���D�z��p�̈V��r��VY������w6��i-:F.�"���@ծ04��!�@e�W��%������*��6��M����3�?���~�z��rC�|�<zws˖.���N�]�}$���X�sCt@�n�@�y��� �����ku���_��]q@�E����!Q��6�k��s¤|�B�*y����~^�R�'�/OmΘK���
u��*�z�I��J��r���F#���>K�|8�b�/�����f�����C>~�dSW�8�ع���N������5�9�:j�_L�l6��RB����k,������[�x͚ۏ��`��9\'ؿ�jT@���ԴM�D�rʄ����^��mM�\�VL�w˖:�59s�'�C,���U\��7�?������ZX��\(��{b�DYT	�^�6��5�=���Xu,���%�ԉ�2)(������ɥ��*�i\4df���'��<<�(4$y,E	O��Ж�@�7A����z>���M��ү�*ӷ�aG31o��z����� �u>P�gh�0A)?�P��<:�'.���'��˻_�vf�� MG?`r�%�ٲ�ܔ�ebL���I�rJz����!�g�_$}M�s$� S�:�u>3��ψ	���<�qo���+�5m��4�{c$,��861��|���)򠸵�g���p����C���Tܾ"��1Q�J��B݋���R�+��װ��C<?�_C� 3���%���է�:�v��I��ݻ��0&���R)_����@�I~3�pN�r��2�n��Q����VR�#B,2�������WZ:M`���g�+j�NtT���p�3??����ۿ�Y�Ͳ�S������(�Rso�h�2��}��x���\��B�%���~�o8ѿ�s�F�o�o0p�8��DP�K�;'ocJ��lҶD�p#à1ݱ����s����5��\tt0a2�hȄ�8��y���eT2�,����A�P.�C8�I&J����j9:j�{�@g[8�����Wg�a��֛@-"gg��.�T��H��a��s�h����,+�,w=i��>��v����� �`�w��{aCn�|�>��!X$��j�R�^_�e~inn>�f?�0�=�Z1���$�[ɸh[6
��jP��@�����S4��):^,��5������T�[�(8f�:&�4:o��ɜ�G�������8��l���������\�j������󆝰�A�L�?U'bu�!�>��H���)-�7J^mo�S�0�n;��8����F������׏�������3���S@�����HS����b���2�r'�V���69�����ʯ����խ��4��,�lI��0�q;����e��,#��v��z�ؚ���U=���VH�1��>�JBӨ�E9"�1���O�1uj��ɛ�^��ĉn:� `v�|di���(|�������'_�o͔� �T�|e�@{�LY)oI=����B͹NN�u���ޒ�������4��w<���������������2�@�I�+!T�������C�w���=���ze�h2#�X��,�F�݅�-���Q�.��D��H�ׯ7��m���7�/��eS�L�,����]��/(��� �|�|�E���+�w�J��������v������P�<���_�]�~�/��s��5��x�7m:i�P�P��\Z~s`�#`��F�N6��c9<�nn0�%�ܑ?�{ak��Q{��_�*:�9���m�X4$e̚�H5��fHf��g�ΘŲ`�U�-�.`�!�v�ɓ�Ց=�����������޵���AB��E������������_�ޟll���)jhh,,����bL�b�X�:����8�u���@�^�e>�-sj_�g�.��cR��:���Z_?��,i|Y:{��?�������6��6~�`P�7W'j��hGZ��
�����;ao����B�_bW�����������v+���������k�p�,fo&��aї9�����%. ?����c[�-m��Fc�;��_�[މ��X;�R�����"�R�~���K���������}mov��v`s�@�J��9��oo��.����9��ʜ�>�"u�B���+�J6!u�+�w+����W�Sȷp>�<�JP��x
[��;�jK���Z���2(���}�$V��S���)��f~��^�n����ɸ���3�=��bQ�^��>�qb�� �bjF۫P D�k�6��kZ�<
ٕ.D�5cvC=�����d�/"�}Y�����[Qɔ8͆88�r�XI���U|&�2�1,�RP�����
�>��i>�#E.��؀���z�ʧM�U�~.��K;)RJ���1����b�ڏ,���qνec\�c���n���P3&�1�Ҝ���\�2�j�%pJb_�u�{M@�ʔ*�������4Y=�<�?��4���y	b��5�������H�<�p�|H�s�|��v��D�wvt��� �j�ϴ�f�� ?�_ҲI`��U,q����﬌R�UN����?�o�s�|"T�C�i�\Y�w	��V�81�n&Bٔ2��5�6��	R��9��Ÿ@����`��G��5��ŵ1`#�d��h�K{Z�fA����V�Dr`ܙ��c�T����OJc����a4�Xm�fƽ�r9��y�*>́+����g�&�g�uǳ���#+i&&YǃqcUs�@��S�\�"U�s���7���&[r�o���@� � p�2�/�ӛZ��������h��/�"��վ�M�ٍ�@�r0y|D�۽r[2Lv-rQP��#G.YQ�������ߺ� "�s���o5c6��~�"A�O��Ȧ�qQ�������tqU�_SJg���PsF]C��I>�k=�2L�D��0��K�'�b+3׃�\�nT������P��-n�7�b����E"[�(2�Rc�K/w�?K���c8L��@�����}4�8�e����3Hz}�+�֭!�� ��Ds�����©;z;��SĠ(f�`�]+WlƎ��H��G0�
T;Rm�hr� �g薉d����0����K0�蘧�$J�:�@4o�bnC��?K0U�FoV���M��@����~�9#M�?��̄Eβ����'|l��M����	w�9����{� ̰���OJN�����$1]�THg�)U
�?7�6p;W6�F����`�+b�g�r�ǭ-aeUȏ����KWg�!Xh*�fy+�&���|���{3ڹ�zΥ�*B6����4*ս���k��'����	�˅��/�BeN�fҿ�ɣ�3�4H�D�Y�| u����$M� �������wk��]����$G`g�����0�(F��Px��p���@n�>TaÖ3�P/��ɡ�d�^���6�����_ƕ�_y���G�3��� r�C��,|ϛ��w	��b8YI�Z
$"Q��'^7�X�s��Cy�	.�,��)ۭ�m�Y�$ޤ���'�(��]v��=��\��?�x�h���b�osSKwR�[z��$�������������Q]��sZ�^�E&�<��=c3E���ʟ�&��~��o+�ZZ�39�[�6r
�tDD�>���oֵvE:�y+bf5����}^}�a������/7g9�ƕA��n|O�|90����r3ʈ"��ϝ�CP�՘��q�3��w�y�F�՗�x9M?��v�6H�O��N���Z^�Ϙ0��*+%�Z�`*��K���P<�C�:�7.�;��lĤ�Y�Om��1�O���ED0�N{=�m,��u��k�7�ρ;��__���
p�#!�t�����Q#�2㖘�C��"{����_���JO�u{�9x�ɤ�a�����W ��5����Cp�Cp������ݗ���K�]���	�o7��^=��������眾�}�)���<-V���C�p�R�0��`3����g@��g�,"��/�H8�����$�J������(���He�Y�nv�"\�8e��,{e�5d{����7�I���
4�n��@�����Z���w�sҺ���_�؄���I�һa��I���5�l@:������?�6����I6�߄O�����.R���7��fbS~-�f`C���do����k%t�DR�0y�f�r���@\H}�N�KB|�rv`n3N.)��gf�q�˰S"�;��?�.Z���#��r?gB��:�.��_���w~�*!Ŗ+^r���l4B�{��0�Q�Bݞ�Ľ��m����gƯ��b��w�|̇3W�Rm�9n�lW>�F�!*�w�&~��}�ڨX����f� ���h�q��?T`�LOǇ�e<[����o7�LW.�����������nñ�*lL�Ӳ�˽��Ł�/	�p6��p`��z&�7����y��k	�E� �A�<�FƟ$�Hї ��(��+��B��B{�!�ş�33A�ӵN/���)���%Z9 � �5���iݘ����R��kU��I!��Uӳ 27-Y�����5��KO���ޚ��\�UV���׋�#�3����J<��3w��Y�+2p�#��%Pr�5�چ!��vKO|�8��֧�6l�;�ZlF�Tr���fI�	[�B&g��!^FW{��d��罐R\s@噬C��뗆Dga�:I)�,j��)	��;'������rw~��+d��g:�(�1�����7l�|?���jo����cc�ǹ/�J����r=�w5�%�N�DW�nȺ�������PY�7(7SGkʡ�l�c���K	a;�!�`S1hw��m�*c�0ºI�J:\i�u$g�x�E�Z� �r2�#^]HwUgQ|:���!e�Z�p�3��q`Rc
�3pV���)^X�рb����f��?f
z���ڎ�5��w��*����8q��u���m��Ib$�niiD; p�]՗���|t� Ff[-ߖ�lX��4����?���CY['���>:��ӵa�@Q�_.�35y���B���g�L�(log���oJ��{�w̨w�$*��ʐ�n�PW4)IV�f�V����_'w[�����m,��V�>�p�l����D���J:R���W���7�B<$v�/b;�>���~���Х}��W���o#���5j�/��N��Q�2\�`Zx�����r �'Ț��AN)4> S۰����YfYa��MRc��t�ZbTV�S�}�h}�a(�e�~ȡ���)����ř?�CU��!a�8��H�,�]��2�֨�����qa�9���K2�D�m�:�t/R3ݛe����"��:m`����
��_-�g���Y$�����Α��bv��R7;>uc��� �7@����U\k�>��ў8���Z�;ߴIh�r�%���A������-?L���;j,/,�V�E�'��ӕܨ2=~��h'+��g�Nl�?l��>�7�ܱ��W�P�DCC��;B�<��r�����4��hDJ���>1_~�5hM�]k`-H�m�΁�	��VS��cI(���	�� ��I�f��W^���)��G�_J���g�ڽy|������� t�z"I���{�����p�����I��t%D+���ҡ����O�}�7�o8���A#iK�6�C���*�\��&���吖����Ď$�����OeC�O���|au��sc�\)�a,OGL����m4_W	9�,�ޥQ����Bj�r}��e�"Q��;(��o-���|+��Z�c�����%��O��YX�Z|?97X�t�a�}�>1u���R�xk~�4�ޔ��)t`�Y}JCy���X4#�k���i��_�Y��0R��e�״�4��Z�!J$/���6�L+��n�:�o6 VB��!�(J�P�Ł��)ѿ�:��ąg�`���Q�"�0��G+Ni�h�zl�S�!�%Ov���5,��ŊC��P*��uo��]�<���!�Ǘ8�V�����6#��]]K����c ���Ku�^�'��ٙ�n������^�R�ꏇ���3�%��E�tv�B�Yr>��Q�Br��
x�`��9ܪd=��JTdHj�/��c�������v��t�P��ׁ�u�۱���!o��eN��--5��V�[zMw��QS����K�w,���I�O�IO��_�W1XN�K��t�^�U�Ώֽ���*�]������L����b#c�����v�fyb��ٟ�2�:�4���f����X�=Z�������@
�,������(#�]��c�^`�zR��`����7���QL8�U\PŷN��!n���O*��Y�>�}H��z�I*��=< �����-?k��$��x�/����]���O���s6�J���L?E���8��
���? ����wƺ�cO�5��gLNB0��,(���	�ׯJ9H'�i�w��0�#�>.�#�%Hn�n����|Oօ����#��啿�/�����~�k�X�>����z�����h�<:r5��ǩ����~�h���+N��+��ǘ�!�qcI�:܉䤏�a�4	����V�4c���C�;�G����y�!���X��y��{g��<���|k�U����A���,����ȞVD��s#��A~�,������>�j/�\��Y���2��OtG�ዧ&�>Gse�{Y�NGe?��e���@	�����Uu���i�LF��v�9.�B +sVY�lR䉅N9����h�!�G?�7H�P�=L8:Y>�^-�ZW�,v��е�8S�I����깛��[�����'Bt���Fi4��כ�U92���f���Rdu�7@!Ô\ta�?�q��G��w8��<9I8ć�ꑰ�l?:IB
�=��΂QX��0�����N)t�����j����27R�-͛0�I�c��;�M����,���s�#y#�R�.�C��&��r����&������c�?]����mѽ&twE)Z�"�(�g�9mCT4P`^��h�5�/����ZM�Z��-��E?'Ӥ�^��%��dt�M��N(�|i�q&=�i�$V�fd8����_��:]�ȉ�},!��hf0Q�	�|/��S�w�ǡ%m� �@	���qxtr�ޝs�J �+Bvu�rc�*����q��[c���6$��EMY���@0�����0����/w[j�y!j�|d�r�2∌�Ƅ��F"K�DQ��_��+S����V�pF\A`��	���D���ջI�T������<`s�ͷ3�B$��w�:*#��O[҉/>�ŪYf)`֏�j�\�T~�1QQ�G�����f��o/�W��+
�p>��[��m�<k����x�L� ���)��␠�^e��C�V�u?��\�k�D��t�pe+�\�����*y0�W�c��3�������"���i�d�R�~�������+�1!ŗ�grY�K�:�BU�Q�Ws��2��G4c�N~S�L5��[��($���+��N��Q��R���m ��x��f/s�;�O\<���h���n����#��� ?���eտ�`�JPs��ԗ�tp~X?�ܰ��,c0��K0��!�� zˀK]��+JĎW�|�b�ss�2o 2ڧ/C^�](.]��Ѭ޹ɢ��ӂW���u�0=��l[��Og��wv^�8���`�Qv�؟���\`��UCzP�Ҍ��r���r�#�k��H3���9����2E��'~k�@W%�SLS�}ZᦑV"`��6ZS�u!��ߠ��*�f=�������~'�
�A�@)�k�F�}��k�{���؋f�}�H^~v��U$�ѺN��D#[A5��5�Q3��C��q��wgt�v��o9u��>��=-E�/Hg9�u���.�bش�fE.�K�!��ŀ|8-b�7�X�9�j}�˖�������"���*�EG�؅�������2L���ˆ���߆"U?�%�����ᬥ4�Q��/��rPR�qq1-�W��I�y��TxY�p�����6⚧#���l�k?��T|�nk����P`�]D�2u{���Y8D�d+a�i&k���F3D��T��'����	��.w���FB0gJ���j�
��2��.��*E��G�\��(o4�*U�z^o�>�Q�����
����O��K��6}�ڳ��9�Dl� �2��󅩹U���0½�4�Vces�5NgY����T�Z�ttML51%\�Q�nRe�KXbᛤD��x�s��'��q7G�,���t��3�ճ� ɋ�=��PB̩Z��Ω]��=՝|��ԭ��T�������Iq���!4ԙ��2d�0c�-'H�w_�M��Kc�wsh��cZA�E3(
�J�)�0J�h}����5�`#8ӑ�M��"�^�|����t�x�ǋ}��b��Qk_?������055�}��}���=��^)��y~�1�jYQ��U�P�r{����KKu:]%>���n"S��ݤ�HN�-|����1ٟB�����ܵ	��gXHG���i�|�<4
�~��u��iA�o׿�2�#���ޞDy)��t���Y��!���62D��?l��o��)�� �Ռl�ܔ�Z9!s �qZY܉�V�|��eL�u���EIw�v���姵�m���� �F�-���X`�ky��+��]UK�_��/} ����o��/��8�gEo�'�vP8��sGt�!�?�I٭^�?>!w�co�ih\v�.������9�����$��#��f�Њ�0 ��%�1'a+�*��]��"��W
����IyM]�I	9���c^�y����EE�J���������33"������~��@R,�,�۝��`��U�jD懗�h֘��9�v(�Ҽ}#?
Ӽ��#�7Uţۥq���z1�5��ֶ|��o@�	���X�ZZF���I�Y�Ʈa3ӈ�غ��o�#� �����J���n|K�O���?m/�X�����y�|��s?�x���;�aҌ8��d�S�ݭ>��Jt���,F8%p�
��=ɟK�aխ�Z����jT��`�n��r�pn��/�κG�΋���qޅ�г���3eBV,��ֻ� ѺWɝ������0c���3�����ď3|���鯛�v�W���Ъ���GCN<X���k��{q�##�4;������}�e9@T-SGI��;��?�V�Q�|���|��og�G �Q����ew���~�=/���X�hx�o�O�lT��N��ۅB��`fј�0��Pղ�Y�=�Z����^9C��t�LߙZA+
k+Ԥ��`�yY�B��[��-.<+`��D>l�e��N�<Rl7ٴ$7�<[�"�O���t�Djc)`$/�'���4I!�%,>~]�Ce;���6�QU���(X��(7��T�\!N`�U_~Q��������3c��W9��!��6���*fI�4�7�>��n��X�����>.�:|��)��������.��W���.n�w�z�|\���`�i
�|ҫ�dA�����0t	^$���_N��l�d����@^ir<�װS�E�(��4�4��9�w����s�_��:(��b"
b6/�_uUF�^\z�珮���[���A��]b	gH�.4}po��ܪ���n�}�k��m������0�5�����s"�:=�N1�6,�Ҿ�`�v�g4�y��yl�N����_!�,�s
���3͖��S�	X�۳�����5�����ι�uo��[���ƥ�՜[�Nn2��.����EV��_��C9�Ɨ��H�D�Z�LL�'o�d��nd��O�_p�w��bS�r��}R�4�7FE�e�{��Sb��ik��6�\k�.��*oC�������
�&�g��������.���N"6�G߃��jy��qk
-��fw�?(��P�� 0(�u5�k��iw�,��D�꯰Q��5<e��I,�Y��6��<z�@�A�LUM-��j{�đņ��൘e�Q^�</��\2�a-E�a_
u�&��0�B_ߏ�@x	*���3ysSy,	#RM����/�`���BKl��+\�t��
��{1�&5[$�z��ye�l�:]���2�vp$�Q�O��0�}��'��б���6Gǽ���~���ʇ����qM�o>P��F-!p�Y�W�H��`�n��'����ΐ�1���6����A0�~�H�I!N�uҨ����
�YQ�򡘜V++���UV�k��շ
�&+����� ��$�[������&��(X���U���Eu��B�IL�O�d���j�PC\XQ�j�I9|��&�l�*L��Z���n��ZN�j������
�rՖ+iH���w�6Y�a��ly�ȹr��A�8*����]���E��h:��K�H$����u��Ch���(-�]��R������D�N:��*QN��s)Rݻ���%�l(x�ߟ)��wvB��A?c�2d�do��u�::��qs�0����Ǭ�~����&�Ƅ�3�n���[0�^�:�_�IN�X/aw���y�#���Wn����f�S.�Jެ�'5�������\f���wG�'��y��q�X��oOM���Q�����,�����N=pE�Br�~�n
]b>b8�i����s~糷G�'o��b��o���^��Ja�&Y�=�k]^̾�{�@�("'��˭z"ڭ��ߚH�Ρ��ɥ�sQV�i�����q'��}�$��[���ף���TD���c�z���}p7�Y4 {BԜ��o�v��~���g�����VJ��W%��jߠg\e�Mx��)�����"�RA��< m���@J�f�A��h ��W�ZXV��(�"|F��F��B�H�9r-AD��
꓁A� �����R�>�vb ��b�(j-=����޴���}yFp��N��d��s��M[%v�ַ72DjPbON��)k�DT����,E�H��=�8^�t���?�R��� eQ.��/�eN��N"f�����2��+���E1��#���'�H轤ω,�*uJ��Y�*b��p��vu�3���Y��Gfꉽw���n�0�[#�8'vs�����}�ý�H�` ��m
l�:�S�W�.o�	ѷg"c^��4�H�D�T�d��ѕ��$��ͷ$��H;�A��������M8�4zH�K��g�m��1 _�u�{�)y$ǜP��q(k�5����l#�V����y����H�́1����V�����@��@�|�&��m�w� �����6�;��m2[0���B�5@nln&~�Ɣt!=:�-�`M�H5��16���ףF�2����]#�hƑ�iu����588���XJ�WN�w�gνʉe{���E���@ �9
�&�\MC	����PCn��r��J�j�B��j���zL�����[�(Ur���)3Wp��R���u;>Q&c(U�(�w�.F"(�{
��.SSTt�9��������^�e��P�O��Ӹs������ޞI<��#B���QZH*�j����$�
8�,öe#L�R�9�%KKP��	|?rJ̈� '�ٮxgN~��p�]�X|O\e�ǹ�p}�j�W�}���:T�QZ�%��uQ�}�(��!-Qq{/����eMǰ&�z�-]�e������8�X�ˌ�|��`�<��(�jf���^$i��#!�����Ʀ7��^�ˮ)���e�:��bBPwwt�	��7�Qv����*0��"0n�&#(L����N1]CbL����bTV�}�f�I0�}�R�0�3܊�P~�EG%��R�:x$UT�G+��ܞ�ɪ%�l�i'X���U+�,�21�Ƒw�ߖ�T�X��L��3��%I���aq�"Վ��UR������͐>:��:�t1��~���k<l�&��.h.0h��,i~��#��N�4�Ir�ΖZy�671J��A6j����H���n�4���և��}���Yjp0t�^:�i�K��&��L㧬��i���Ox̪Rh�Q �.�.|6(> W�p��hG���=C��#����@mx�5'I��>ё���9�a����ݟz���q����Y@$��p����چԣ$5��1�z�z�}#n>��i�@UC&W�RQJ`� ��#�E8�����&!���	��������	�.Q�qr
�z�{�������L7�}�?�ǂ�@@�9X
�����s�h��JgՏV��X�����M�'�#�'�9{��ju֚C�!I,,[�{s2P������Ć�U�X�̉��+���
���Oϕ/wRP�����Q�_��*8S�BS�U��b���P86��� w���$��'Ȍ{�c7����⪨XQHu��7�o����C,������J8�ǔ��?���VG5ے����0�LM���}D�?#R[k�A�'�-ނ��E�����G��72ӥQ�̇�?���Jl
cj�i�ƨ��m=����8�q��@'�[���~v��	6��n����C��p���$�ؔ��|���ӣ�����] -��ڊĞ;ؖ��l���.�HtCҸ<R�4Wa=4@*_P��Fm�Q��v&��SK�I$�zg�P^�n"����m��r <�h�"v���/�`KwBũ�ՌTfw-��wҊ)�~�߼��W+���$�+cq��ޑ|������;~����g�{��}]3۬�#h�'��w��s{���)�����8 #�R�
�t�WW��vQ9�x�¤)`��$v�mL8�{g�$![��{� X墲)�QTS�9�~��צ�`����T�lgDϏ���AF�0��
ط���k��c6�{���`�����������/���.|9J�4�r���Fb�I�Me�%:���0����r#�])��������F�{V�����âGӭ�5�V��;hk9Y��hnۦ��E��!�g�,��>�o�2��Fʯ�G�>k�:�t��Nnմ�L�[P�]��3ɸ���a�p��߮Tօ�$�q� ճh?��+i8ڟ(����$PL��G�_{�^�i2~���(��G��Hw1��S��ف�M��6�G$T����b��#$ 0�n>�+͒Z�c�:aݺߚZ�+�{�(D�u��|U��YF$HO��TEQGR�.kE*�+n�f
ڟ�t�;]��h���,ڡG!�3�\�.����dn���;�<�֫	�:�'��}q��߼<a	�Ka AQq}5|�&ܰ)M��H��DݻS[A� �:���Y塕&�/���̀�o�������?�Z#�W�ۍ���|�����eO���?�$r�M:m���"R[;I���0Y�\�B'��$9Am"Q�m�'h",fԥLA�:��D�δ
e�/��� ٌ���.g;�T�q%W�OU'�O}�8��.�c�yn�����/�13y6B��CU�Xi5��#m ^�@� ��㶄����O(����J|�iWL�c�ۦ������������p����w��Nz���1�K�����E=��}jJ�ǳI+�f�P=F��ix{j�n��
��*��~V�KFІ���Z��뿺�c 7����^"(y�0�r}g�UGz`�����Nvu%�x.��a�����p{���6�>8:2>�~����8n԰��ķ�����g�5��! p���������v��Sk�z�/_AӦ�(znQ�� ��t,؄Mx�ݧV]��p��K����p�_��qҍUT�7��Fj��0XF7 lߓo]��r(�3Y_ޝ¹�n�l�(�o��چ��]�@�2Z���({rf`�2ع�[^|�'����O�וE�a7�c�K��k���@NzX�6Y��9_Z��!ߛ�:�ڙ��W�hy�$Í�y<�5������Q,������k�H��}I����DD��b������k�u�'_%$�S��P-!�G�] �WJ��~I�c�/���1=T�C���8�J�s�dℭԞҠ�v,W��<����Ϫ��e�����w���:��ᄢM�˗����s�rKI��C��Q����'	C�C�s[Z��AUϡp�Sx�S��Vh���!�.�:΃��:���-�8+�o����#�Je|�P���dl��ZH��m��� 3/�0�����m͏��y`�G�`�iz�!�KA����P�����<��"qC
��q�تP�6�'�8O.6+�t����]S��UI��XX�Γ�ڛLd.,'
j�j���E�R�t|���xN��kB7Fq������MQJ���dI�Cgc����~��k����o[5���AA��sZ�u��)���O�9�$J��P���A;��1��Tp��B&���0ݳݤ4��"�k��2�+(�&�2��Pc=�����A�	�wn������F�U��O���.YƳi��#�r(��/j�o/��r�6Y}6�Iμ�	�n����a�U�Sл��B��╨�&:�`�	 ��<kF�?ooo� (��d�J�<�lo`B�6���󆤽����g��"4<>ٰ���7���B�ͯ�v_�[-�F�|��u11s�Y�6N���B_�ⲇ������Kl&v��ˏO��F�/+0#����a�/��M��]�.6πgK1�`f�+������t��0f?�)��W���Ĝ��~+T���}k�ة��8�jB�`��2���9�N�Є<d��z�s��}�Q~+:u�5J�d���5�����-��r/�ۅJ1�\�[��0�*{>�_�M�������5�=|�i����~1���af�Br�(kX��̍��E��oѦO 8��Å���P�����Bm��(�������X�1�����������b�Ht��9�iE�\���:|�T6L-7R��_��^�,ry ��*��Y�����b���u�Щ4`n+���6j|�t5�ͦ>�6;���bz����������{m��Q&��H�z�7
8��bed������u��ԁ��l¥Kܥ^Tҷ�5�����(���	bB%�$�
�,j�3�z%v��Ln��:@���??�б��ڡ
�yP��)�ev{REG�T��a�]l`�`4�7�PzƋ�#��ԏ:�~h���df��w��~��S=	x��#�g�"ؘȖuH(#�c�P�q/�����@��3�	�c3� �q���gX|���%�6kZ�����Q��0������&	�����<dt�}t���y}�~ˆe�uy�Y�C�8]
�SΤ���_R���w8v�?!�(^�]Z5S�8V$�������[��q����!�@��Awjv9�(񕏦>R\r�P%��\�[8�mA��I*��У��K�A^_��+3�^����W���|쭟-��&x����z>��)�ŀ2�@���v!0 N����5�������C�[��J�Ou�:�o���H5���X8�Y2�'��]�L��~�{����j�Q�T)	�7����:�jXQe�K���YF�����m�+�kV�z~���tQ"2o��?�M5w��Z�.���~̞�{�H����ݎ^p�	�͇�>�$z߃���f�̓������<�@)s�/ vv�����B��8V]7������Vԯ<��D%�CA���%���X1�9�c(�՘����e�o��eLI�AnV �oʫ;4�G�.�?�Mn;�9�*�R��#�=何=<#�"�?>qpSȰ˫�j��(� &lr橡v#^�RW�]�����b�����Vح�Q��� 9d�A�����R���)6`m����Z��%kب��,
T	š��LT�(�KaCp�|�Ҵw�)t��;1�J:U�8�0<�S�R_��J�aD��o���q���:��U���)��#�4�Л#�E����E�x.��,%8u�S��7K��|�N�6fS��u\}�Ex��K�2h�ҳ��<܍%�=v�p���lli<W��u�p�
[h�"���+-a�;[%�������G�:�8
�~�n2R݋���T�Aq6�=���ȃ�?�I�|��믏�	�Y�:��%��!�fk����c�?�֐&�cf�-�5�-U%��1�d�iF�����fW�k��(�������\Y<���N(/g�[������'��W��; ����ּX����v��W��o%���<�yo��]g�V����R�Po��att��M;8 ��qEW��>h؆���r�����2m3w���C�zg9k�$U��.��6�R�f�`���~1c�E9ǌ��F��V��qKt�#j��iK�N&��Al�h��(��,��Bʝ'��^@��#�B�&&�o�?��W��jQ;D-]���8 ��N�iZԢ�w���Q�`�Fq�^Ծ����]<��3�S�����r
l�(����4f�i)��&+w���@��
2&5 m����)Rp�k+Lc|��(q�O���-B0�$����F��D�p��~^E	������x��|z��(�$db����r�F��AL�Zh������`E�v�`��.l�=*�ָ�ᐠcg�c�4��z�E4#/y�[��e��1�0cӲ}oH
�'g������N$a�p7Ζc.!�P0y��D:nѷ�SI�*j��-�G���n���|SbZ�iV�8a��P����9�CS��*rH]�~N'�>e��Nc���)�$� �`A��05��w��3�*+a�@�+̣e9�Tޓ����ͷ��8|Z�pc� ���6~�W�(�0����U碩Gg��[�875�G�c���d�8�d4��{�>���܀N�\z��a%dd�Z���~���U��$���M�_@�u�~9So]oS��7�xXS�9�8�+��~���&���zp�w����Q�TK�����Y"HN����jI=��0�e�$�P�5��U�⽙�d숾R3`'�.k��~ �����d�b�����隍-���)	{R1S��D�x��^�%&�vf3���QBN�mHD��f�HB�߲�f����b�~�1^ �abbG��@x��l��r8xAB'
k+�?{�jR��<4�R�]�zR�i������0r��F�r�ǡL�f2h.�c�A�e{HF���o�F�ϥ�=7�q�g`���H#X�hG~��0D0qC(�f_x���Cu�H����-��*D�w�D`�ٰ&���,$�@d)�7m�j�5�l�kE�4f?������Jx���{?��Sw�y{����G��s/:��2�FDA�
U�9O�}�ĩQed�~"60n���IB��cq�'o��i	SR�S���'C~������/��� '"��� O��}�CIP�Ƃg}������p�5�=ݝ:���ה��%$�H	H�=��>+�����鉌<�i���A'8�0xi��A*TT��H�g�gl��i٩������D����}�ȯ2�o��{A��+Z$0K��� <�N`����;�hӷ�K�i�Q%�)�X�v?�O�D����6�k�	�����#��w��js�
�����ӆ���a��;#=��8u�r�Ʀ��7���ɸ��5	�%�X)�	ײ��`Z��;q�RI@j�.Z����,�����y��t��}E�����|"�u(��39�>.�����&��0�X~�IX��:^����\E���E���_nnn�
rK��h��Y7�&�3f�c�����DLcV.��!�`�h6�>��h�4����?���\���v�����Y�.(hv��3	Y�0�)M,g��L�_�Z3��B��8��Uܷ<�3�+(�3^^��������:�}%�~#�n� �K|�a�gэ�@I:�T��vgSֳ���t�D����w=J���R�'X\1v��l����_�u�Ng��Cʮ�̏��}z��;(���o���7�vҶZ�� ��9���h�S�z���/p���	�gfʯvZ �f
��뻦&������=�ôQ�·��-킟y�	-N���'��}�1_����z�/��}�_�'�w0�Z��b86GGF������0��n�d���4�?��4k����k=�;XY���������8bm��0l":�ݭ���X�)�ל��-��22];�z7Fw3I�������PͬϨ
����B��G�Ui�ǩ��Y��	��F�%�K��0>�M�Z�`/�?ru���y�����Z�z����N?�f�.r��܅!J�-�5�{�Xx�[��,�G36"�|��	~~�/��6��_�xx?��W##��sarS�������$D�����2�-�]6k"P(#�f�m��[�����0�=0��{���$����R�t��&&�>���։�H ���bu���i{?ʫ�Ӥ����l�3:ZI9鵠;�z�C4����~���Qs��.�&���@��Q�l�H.�yHC��%��& D/���	��P�?���:9 ����\Y�+˜6}oɡ�j�hZ@5	���m����J�# �{��?��wJ��%2,��#(��"\.��?�>��!��]�Gт2�f
M4���%q�H£�1qˤv�U,�&d�oiP�B���Z�Y���㛀�� �����>���tY��Of��q���>55���b�� 0�P|Yh|>�@?��\�j#R�_�L�7k��W>�J�8޴R+�w����+�{xNi�xB�JaL/>|�Io5��H2vz)U����MO�P�/6�7?g�Z��� �p��p�j���)V!	Rd fFp��?����w�����2v9�mD��D`EgǚP�^|�`''�+�\�N�x�٤���~H��n�C�*���q|_sy����VFFO���v������ب%.�rFLө莽]P`z��+��M:�Ɋ�˱�P���٬������]m����6���YN,nU*X�x�ؽ��]+�(�C΀���/��~��̂�k�ݣ1���cvn��!�FQ�e���`P]��C����5A�䈓�OӦ��(���(֧VcJ�>�
��nm�esA�Q�͍rt�ŵ��	�{ew�ljW�s�<��E�G��O������EyF27���j�v�b����
���	�EL���z^_��0vG3�������~�)Dk�T*�i1FF|�K����`�01��3�Z-��4�$4�3��x���W,�l�� �V����a�g�'g;RhE�5V���뫒 y�&������*���J�g��W�y=*����X(��Oo��G���X{a!J�ƹ�F������-0�Pnl�]p�9G�r�qc���&Q�[�������p�/vHG��@ο:��zN;`s\�R$��`f&(������U��	G�|������A�����sk�dH�T�Yѳ��h����l�B'R��͖�im`2��`_\'��ʊ1��˭䀱�fŠY�>l�����ߔ���F�����(�˔1������S�#H��ͤ*T�Ȼ ����d�j~N�����S ZkX�!?'t� �[U14Lh�]413�������7z��B�X�;����X?7�����&��z��Bm.2�Wr�[�.ΒV���zz��>�@W*�G��w��g"6M�r�a�i� �e�����7e��L�Bn��D���ʩֱ|��P��:q%���щ�N1�T���q���E�)~9/��o5�pm�p�Ϟ@�%���"N�+��8�a_��^���~u���Ѻ�S.kE�x��経� �h��Q�[W���U��ce$���m#*}��ߗ����`�-��%�"m��[s=���!<�b�[�OY9�E�R�!� ,s��  bH܀��!2�1��g�������jx��a��5r�1D_5��S���j��ìL\\܍x���m������әx�7��>_����][54����gE�o�7I�5�ꉢ�Z� /k
�a=Ůڰ$?J�{�(]��&� Hz���t�Ő��*ä�KC?�'B�����(b�DjL��'��!"iS��Ϥ�'*��3�2��X�U�@�Pbc�%t�u�)�Kw#�`N���IM�ZX]���˫|y�8��9[Qx�Ho�<\���P�sڐ�1C���������f���Q��Kp��� =�/r�v�A��,�Sڑ�!w�������|Y3v�f[ږ
��rX�\�h-�S8ևs�rD:9 ;����([]����hl3��̡�����nM�p�x�zo�v>����j#�R�W]�)m9��Db��	�sN��蕚��Q<�0.&6�GN�Ȳ�Ϥ�����Y*�
fh��DkcK�y	GG6�]�999�2�1X����G�~��L��+��Zt�������щ ���I.GGG� �f�7bC�t���*D�xޤ��L���/*���dѴ���<=���BCa"8|�ӂJ��YHt����5��x���O�e>w����lcp����)b�Fp�DKf�~D|db�4P�쓍�?7��4A���P�B&�~�#a�^�q�,@��䢊�f8 \`nn���ڽ��@ӎ�U;Y�E��6׫�b���h��%�hj��Gg0��__�X9-�Z�����kT8=_����I<�j��n[�a�����>E����lQ2��h���lV��H�=���Ÿ�]	\F�p0���G��=\;�Tت^T Y����r���ݯ���&�1@�K�����}���#��]�6��&|3�]4��2q�l�k`�FE���s�yH�&\��,��:�hli�l���m��!�-���ڮa��-!��Hw�� ��t#���ҍ�]��i��Mw~��z��C��Pֹ��sE���5�F�33��R�^�&�!�ٜ���o]��*B����I���V�B�u)��d^A%z���f���Jk�D��ν�SY��B�Td�r k��쎑Q�bx*��2��`��Z��v��8��_��BY�Թ���Z�p�2_K�=���{����G���d�o+��\����a*HK��zg˾VYLѴ�nD��3�
���'��=9����oo�oDJ��y�ϳ��}Lҳ���s�YAMB��[W���4l��ݶ�(�0?����W��%f�W �"''��X�����`<4d�勥ا�Թ@��Wʋ�s�����	ּmq��Q���*�G���ŶE9�[�{0�V���_�E!�y�YD�R�A���*�J;��m��rm^)5���H��ތXd*���]}Z�ԑ�9�/}ߗ��a==33���p��Mt6�Xaަ��6��?3�U6� ����$�-Sհ�*��KE����'撴�#N!Kb�gL��j����M���0�đ�m�ȋ��Ig���#W�@��nP�'��A��q�ۙSd�;݀Á5y�X��R�f����~���|I����=��$C���_9qJ����hMԼ���d�Ywi���84$�x��'6��I~{��"M���)��d3RR�ْF���%�����Ȗr���@���a�g�?�LP^|�%����K2�����K*#ww���Q���xm���U��p��p$;��Sp�z?|c�K�|_�^�d}}Q�Y��F��2���nw���R�Pa���a�/�K"ڽ'�]�5[_����>���uCT%[F�F�ݿ���f���3�i�|���F�����&?ur(HduY���2-��X&���(,����'�C'���Hl���O��W��I�-���(E=<��AUm\BWxF+,5\��b�
�[��)�FL����uk�͇�����9Q�2������5�s5��5�:5&��'�ĒVlT9��l�/p6\0��ب�Ă���(j-�1�-��c`��Ы��y�V��;&O`���[Q�r6��M�NQh�������*���@]����j�)�J�J\�����fx�_-(�Ωm���:p��[��Nn֮��e�^ł��;�}E���]�ll5�pr�`Mm�Q�Ɲ4K����vO�Q��a��=����Op��}tq�\��%R�?4-�2��f�7�*�����b[!zhhG%�7\�8�62ߓ���L����q��:OA�����ֱ֮2�v��훹�P��(��r`�}	5�7���<I��BC�l���9�Ρ
�e��zS�E{H�\^K�Ͳ+٣��!3��aһ{Y �s��QQW���mK���9*֨���)Tb��0�{���!NsɆG�T�?��Y���$êx�-N�
��À�NHKcH�j+VN?R=�o���B�Z���ұ�鸿�\~6{#vP�o��4B�#~�+ڽ�/�ʔ�T�?-��*#����{��?b/����+%����Mvӌc`Sly�Dh���xr~>��p�gY4VvX�l������A����D��"�O����������s����
CKY�|":4�N)k5���aq�ט�v�0�R���i�_�p��z{(����°������T*��h�C���:�ۿ-Ҹ�9�x]�ǂ�1�,��_�w�{�:(�Jٯ���W1�TC��AE�܉��l��!VA���0��yo�����SR<k�����P}��d�o/!��u�H +=��r�5�Hݤj���V�|c�j��dD=Z��{��^�����K��G���S�~f馾,#LG��G�|CCJZ�1�"]�G����h=�W�����(����?�����Wl�����Y��q��8����%���$4u&��eml�>��^z��G��|��$W},���:}���ձ�9�zODA���>R��'��x��&�a�� y�0���-��}W�+�p��x��Y
�Yq�ڙ�	k��8�2{s�'�T�P;/�����ϖ<����7bF���5�Ι�fPU�wQ�g-��0���1$�u�gR(�-v���F���{sYD��U��6�hʓ�Uu9!��6lE�䲚 7�H�O�2�����[x�k�jDP����'f�������r�
�mw`�y5C�:�9�R��'K����L���
c=�\��R�O��n��N���^�&z�����7J�t�Г`�A�"�dq)|�o�Y�\M��Yt	XM�A����1ٜi��Q'otDvw�P��ʈ_Ζu#�y�.l�A���?t��!-�	d����"����KP*����w)�㜬��0�����``@�Z���5��_҅���S��Ư��ğ�\LX��H����+HR�b��
	�yA=V�XAH��pz���'������h���2�C �������L[���$*�Ac��B�Tє��J����ug4�l�(v}���y�D����1�T{����{�)��W+�����(����v�o�9j�ϖ;�����ch�`T\���.����Q�y��e~$'eP�Z���瞺�����w�bY�Q:S���
\�v%�T�sRW��g�^��GO�
 �3��Ⱦ�/��^��{dU4�#���g�z�ՈL|"qB[�7�^u�'17x�ј�dC�(]���c�cX���Th�R^���nF�v�rN)��6�q�����͝���Y�$|ߒ*o�`L����>���
X�~����j�5�	u��i�N���HY]p8�I9��?.��®�AA����k��H�P1��
��Ȁ���m˛����o��!�����h��)��tI�Ĳ"��E�6x����W��0�����G��EF����Ʌ�����s��%RQ�)!vW�&���:��-R��I�K*\�)��b�leM���sz�B�f(��,/�ײ� &�z���]��b����n؁/�l����մ|0��ڴϚ;�j�C��:����:���|�
#5�nh�������gZ�E��bU��$,��%�q4�+��F�/^�Ew ��|�B��4���uW��(�ę�ۧ��u���F�3dK|���oc7�/[$]�w���Fg�w!�v(D/�'�o�嵇��(۪+	[��$-CD�W��4]X>Y�h"v*♓;|uV�<�%��-�,�W�iJvv�5�)*��V��7�Q��'"� e) ӱn���tt���t(��ө� rc�Yϥ�����1�D7�ĉz k��v0�w{89�d������2����	+�$%�co��w1��WW,|=�����#�a�kL	
�Z�͉��@�._"xd{e�y��G߾)2�|��􇨼��Ak�c�gA~Hg0�nXs3?PjGBBB��%ةz������p�f�K������a������E>�z���\���Ѥ3�������G�)���3{nͥk��Hz{��TipDD���èV�o�l�x�`�&�M:�e�F6�u����)��Ed7��0����\#9E�X̔L�Gm�)Z]�N��3n=<*���m�1^|�U>�I��f�G�0��V�����~�}gTI6ߩ���}��ۚ��\61��<�=|=�H�0r�I��p5�2�6#FD�k���R�'͍ĵ��ROBBH������g��P��T��{?������%�GW��G�@�%/����8~�'�'ˣ0^��C����~����D���*��I��1q2��(ގ`�:��r���|i�LD��쫃���n͉V=GA>ը]~T�p�͖�dȸ47�E���� ��2�2�!8����!q������Kt�J�Ԁ�mKo�Y�*��|�O+E�`9W��yҊ@o����\䊍	���?2TeO�ДU��b��I�<���Qu�r�`
�]w��i�$��g���F|���ϔ��>E���WF���	��~�DQΤWXlPN�5
Y�A`�N�������Sa�� d��!��kj|�=n��ӻ1�|>l*�t;��H�9�1�pg#�4�r��'���ZHb�ecTmЭ�-�����M�,Z��ap\E���>�$K�~+Y��ѫ��'>(�񉶥�������I��r��L�.���$m��+��{��cΠ��ǝ6�J�����}��F�������v�N#�wz��/*%"���Y��1XIOOҬK�X��`�C�ݧ2�i4���:!���[n����h�	�؃ϒW�N��r�M�B�0ޣ�]%չ��p�`�|����8q<c�/[�P�_��ưP��~��7�u�A�#���q߃&ei�^�%?�@i��FN���������F8-�!uXS��<o_�#�>�]�cQ�E�r��������aHL�~���>_�
<������ W/��pԨ�h˴y� i�lon������꾫�Vv%�IҸR9i>�bF��G,�eפ����XE�S�������MJM[��6��%�����ֵ�X���>&sO���������3wJ������Z
����K����O��0�/TG��	Жؕ�R�D!�1+?M� M�QP}-�����,{���;<�f6�1�|Ԣ�2��C5���s���ۓ��÷�K�Bi�(*wͼ>2�_�����&8p�ս���ۨ��r��~�) svv�Ȫv뱔S㨫��΅6~�=l1�C��2��cͩ��`�vr����4��I[�Nx%���=@m�df�T�nhP��u�]��g�@z9ɵC�Rbe\��w�>�ٶ�?C)�m>X:H<�o�5c��ÌW�����ۂ��c�7���F����Gd	{�:� ��qy`x\�Ƈ�����yf�l��}s�x�{�lڥ}�}�}su�Q��KE��;�����+��������Du���f4�B�ѣ)��_M:ϩSK�2��F6s����p�dd۠Ў!��v���o�7~�H@��Gr�^�O/k��W�%L�~s��ߞ���WE�;��}_��ƴ �[W����+0�:K%4B�X6^�f�{�����#Ô	6nV%�W|}@�o�;Ψe��/#/�a���l�VE5����\���j�i��3OG�;���\6��S���j.2��u�_�/�����w��@�i�n�*Wc;��S�B��[E�X�����vwBlvw)��#&�Q�%��l���{��3{~��;�vE��۟УRNm��l��t���τ�~6,�~]c�{yA�5���؝�3���}3�՝���>����d��|�G�-
�! ��']sܪ�&��@!Ш*+��V�8����e��7vk�A�+$��F��&�H��<�mݠ�hE�W'��P	�n��ݻ˔�}UX�"�t����8�E�-���B5�M����O���g�@O_N�(P6��C�CyʥDX�y�^���
���v��!"u ����9��MOOM߷7�/7?P��G27f�F �p��Up@�sj��b���FB�h��.kEhܹ���dx;�t7<�4�����w6˞��Q��{.��Ĉ19����|\�:��E&��DL����>�=�S�p9�X3�+���8�1�ڍ���<ߞ�	~C��+D��֗�pz�$���x����ߎz�[��ټ�A:k�� pg{#��(o��6�E�CPUd��,�i`�u
zS*W��4v��_���˂���MT�&gf�ّ��X�9�3j�d�>�ܝ��l����%��	�Gy���x�6xG���혁O�q�u�ȫ[84�	�rrJ:q��Q��x@f��d�����	�$Wn����%ڎ)����S�^'�n��L��-+���:�)3�idE�!)˺n}Xn�4cM��4��di���)�	����.��� �-�ק��lv���^)�ڰ�_��$ �/�)]ۚ���VP ՐׅT�}���n0~ty5?�a�F�vye)��A&�o����N0Eq?�omoǡ| q�M��jXv!�fi�Aɟ��/��z7��&�~p����V5L���-�Fa}	�o���bɋ��18��S'�P�������k�׬��d`��*��I,�u$��<έ�]����e+��J���7�3k��J<��%r��X���p����$�e�⽢Z�6!ɉn9쬶��4]P�b�������7�h\V��q|��·=�D������x��y�ײ���;J@%�С�᭠�,ٸ���ڄN�c����9���țm�/��������N�i&w�i���`���gՖ�y��@��ƛ��á��?8��(�o5V�\5ҩI;%#㳇!��3���GF���}L<�a�q�G!��pE�'������,�D�%�I�z3Zw�hE���X�c#������0���l���#�D�:��BK3L|��!�DR��*|i*����71|��� i�VZ?�'S�Ղ�/V���� t��Y��E�ƚ��#���j$��$�V��2G��~�(g�����-�hU���Ig��������إ�C���_�)6G������o���+�-��p0��xYUx	�x�����XZk�U4@i�ڙvd�6z1�4Q�Y�����#ƐI�~���)9����o!ʭ���.)K�#4��%�_��
�w�H�/�P�,��@n�*���9������,�q������4\ ���S�©����k<x9+IˀґC���3jk���� ����pr�7��g��y�a���ݥ�o�g0�q Gd���u[Kl��*��8�,�q蔑�Q�T��ˍ\"��I;$�H���s���-A����@Ә�!��j�&��5`E���E�D�����_�)%ipp�F�!"0}"E|�3. �V����rp~_3p�C��TE%26e;[��7K����y�ڛw7IocW������C ��~v��J#V���_�W������YBV6~r�k������+����(�&K$#��-R��jNY[�pb)�r(� *�e���C^�zݲB��.�O��-T�::$ ��:������>�3�eYx�6xW��eV�������^�M:��MD��1Mp��e�7�;o/�@S�na74v%D��9����D��x*�P�L�S���l���S�~u3^M�1��Q���Կ)Q���v������sO��-��w��
�t�U[}�5�������:�kX�z#���s�{�&yj$����4b��b��ܴz�%��4�K�B�@�-Eķ���Zr�@KQ���҆��RD����N� U�y�e����z��]������}q�K=�DZ.?/9�VV�z��X&�~9�vۋ����@���0����-��^ �D��P������ɷ@O::Y��~b� �Έ<���oH�\M��HYk�� E�>w�z�"w�·k���LG.�LDL�Z>飦Me����,��|�~�!�5�a��2�- ^�o�ݿ)������������L�t�p-]�m�v��!�Bs*~x���O�PQl��CG�J(Mm�&�\��\�[���`}īt{C��	�;&�0R|�bWO����c0�htwk�PZ�T�\��P�P4��L���ח{q��'��z�њD�{��9hEXI���d��a�ex;��WM�5�`�̖�6�t�_so�j�[����H`T����ͺX�F����k)w�e>����tpѤ΄�(O�����+��]��ȴS�s$v��{�^�q+��uw�x�F�M:2R�"���S���k9x���Ǡ�z�c���%���5E�s�M����}D�n34������`$^U�4��1�(�P_��k�M/��b���!-���w'Xˢ���1�3Y�aĨf�<�p�d���c2Ǝ���"�e�`F�eI�i;��~��h7s$~��ar����e	2��I �55��v�^ <:5�:K�갔-��'AC��--r��D���
 51$� � �{�F˝��ů���s�z���t)Vn]\�����}fk��o��/pm3��VV�i܊��t;3\r��JP�W��u�dϧ���@C�԰�5r9�QNi��Z}r�k�r2��9����[���i�ZH���Ϻ�9~�n�c���c3	azϓ��B�-3og�������+�j�����>�}��g3�(�n�KoC=���ݴ�kn�a�z���V��%�w���5��|;�&����僋�$c��z�!��e�TOc�����7���G.�_Omu~���mm���B����"\�����T����-�WF`5ޤ��Q�=.���D2�~C{c�.�;���:��b�PJ�iE�g�C.�.��;�J�K<�|A��Sf|�To ��!9
r���S�A/��tI<&s�V���&���ӱ��B6]���="�g�J��<�@�iL6�iy`��M��
~m�"<,�V��f��Ygm ������M�����z`&g:
��$�����?�C����rc��ܓl���y��y�V�4�C��x^��m�|��h��1�sR���*!Uo��I5�kj" ����W_zy�	�
���v7�b�>�=�/�Du���+����T���ۿ���Ҭ��)���]����,���i�[)�_dQ�+� Z�T��ifό���ܖ�XE�����T��k,�c�ǿ�������?,k���F��C��_�5 K*���4�ˌ�RG�3.b�H2�S& X������o��
G���`a�*����0@��x˿���!�����������-�2���?�M�7S,Ny���#��춏�R��r<O���ߕ䬚���p���n�g�PR�j?"�d��v�z����HcŽ�QAR�[<�}x[�|��: Q��ܻ��x[9�Y
p%e��(�%�l�8.�G�9�0b���MQ�N�r�o�>{��D�JmLczY1��'�> ��+�7:�>��4�v˰�B���x��N7X:�I(�q���`�K�\0֏�I'�绺bخ�#���?���%n+vǏ4a�.��fS��U���?�mT�iE�$a�8�47�������N����F��;����ᴯL����Y2���߸#`��
�w_p�>>�?+���x1!��������u�l�n�3!�"46#�x*jWFW�~����X�Ku��k�1��qͿ�k��LhQ��nN6ޡ����z����a��k����P�Yo�$�I�ysZ8>8	;��o���e�ܤ�ږs�)�s�W)M�`3n��^!��	�Zi��sc���3�av}�r�k*��+H�wk[,�b[?x�6��p6�*��
E/4�����:D#�A�K������q��[-��P�n�����"P��G�����,��(Dͫ��Ȟ�i_��R�W�i֦�2���E�XD}Ʋ~��D�F6�\h���2�n<f�ޞ�9MSɪ[idj�yE�+1�N����!I��>�x��G�e��*�;���k����gQii�(�j4~�|��Ag_Q�?[.fs���a��ĳ&28�U�f�ኛOK�5?��Io�vv��R�E��o^�h)��/��d�{�k冚>�U�����63@#�1�}>J�4�/?�WS���ͮ]+�/��\���x{t�S�s�$�yB��s��"ݯau�s@��l�W6NN��n��m�⾛_�«r1H*QLp0��ba��;�z�?-�o���ƯO�f���-���?���ډ�5�hoy�9%����V{w�#"O۫�q��A*2($�c�1I�rWv�w�x�������{3V$��k�H_���_�T��?z��=ݘ�I�@2
��;�����>���&�LSSfo��i���Jo1j�#����P��S�Y�w*�����|x�'�h�+�/�+�R��~�[f_�;-��-Ҏ���������ƕ2I]��~~#m�i��v�nk%�د�m�����e����g ���fY��d�Ļپ>2����r��5K�����[.������~�%	#
)zZ�fZ{5�b�T^��V֖b��pH ���oȼ��D�X�oF�T��jxЉ!p2�^��k9ra3E���^�4Y�~2��`��{p���إ%mm�e���?��	�f������#h��f��g�~d5�Ȗ�LϏ�r՗L�����)2�N�)��񜭞�E`aD����m~�c�;�z�?�v��jf�ǝԩP�G��cW}��JƬs���dt��7*�7��`���w�J\���x�)���~N��ӓ�����M箉������˩E���GZ�>FFT �6Z�ݮ��_y�GGz�2I��f���!��� %w�b�Q�P��7pU����d��&Q�&n���`2��O@f��p�e����DC��D�5���OD�g�1�����+��SV�GG��.����8�A,��	�ۋ��[��zӫ#�:NF�RQGGGe8����:n������}�ߜ��?����e�����H���mhÜ@�[�N�_�n%�ޝ?X��NtS��D*�ȸ��o T\����� �o�Ji;�R'VUS3u��l��Wb?
b�OJ3��&~���z�L%���/f'-�0�_F��!_^7n��!�t����R.?�/�$y�fȹ=�~]�.M��U�G�SD!�أ��M;v%?��*��J �Q�QS� ��5\d��H$��]�}�:�%�?�y��-�<@x��s���c�؁��B��3j͏m���\���Z	ږʟ���l⵬k��H|�L�%�c��x�5A��}h�������ʉ:]�J��s
z�p�D~<ͺ��e��M[��:��BEaC_��Q@���P)�&���w��y���%��1��DKS��,E(��h�&���_X�{:�-y�!A����tkcD��b*��"plL~��c��Z�7�.+0���.���Bb<�Wyu��7�A�qAI?���_?���|�c$H�h�x�]��~���l�xX�Q�����B��~��Y�,� V��6�#͏^Sc��%���/�ZC���J˅��j���=��TE�(ޑ"-��z*H��,b�����y���Mz�����e�b6.H�ңdcL�^HKj²F�L�5��ƃ�]/��[M���o�O⪿7�K��9���f�X|������t)Ywi�^"}S��,��"d�uq���t��a!�Ґ�b�\i��&�M�?i��B�ܼ�m	z�Y��ۼe����!�:4�ϴ���^�d+wji�Hf����.���x:�.�tE|���-9����l^������{�v����� �����?5H~~z�^�+���?��k/��`��y��vC<�s������C�6KWVQi�1������G���J�&��h�L:ބK����-�-��I�zL�w2=��D7�/��� mtnW3��P�P3�	���7hhhvw����:ff� Uv�LP��"�25bb�q*jQˀ��V�jОF�k=���4w��~a�~���;$��+�W�aN�\�)��Ĝ|~�&�m��7Vz=���I���K;v�W�o��
7qi��Ŀ�{�͙qE��>/D���af�j�l��Z.��_����T^Pm��37`�P{C��}�������FI%T�L�m�����l�䵶v���Ա��Bc�hĎ�~`����*��@L����6�QQ��!��3H��\���5��S�P�԰l�spx��v�� ��Ll�X"���p�Im�&��������8e�	7t����v�ł�e�:�"��@������́� ���P�.��!�*�q�`yc/�Γߩ� z��A���K�B��t]��7/O���n��O��2�)�%uL��V���.R:���F"ΐ̿���|'KqS9C_�H��6Oϑz����C�J�㢉���:�o�[=������\N����a���n��k�%ԊB�r��ףݐ���o�f�v`]�$�u��Y��$�F���I� �#��H���XG��<�)5��y�@�v?�mҹ��D
�N����3���B�*�����dϧ�-�-�1ҧ3�z��9~VV��mQTU5.��q�R3Z�ˢ��UK�Q9qqT���Γ�y��V�>�k�-3k�[��1�;��n��f�g=/p��[�^m��TM
��,YO�����0k-�uE{�Q'+���@F1���ɬ]�'s�����Q(�F��`�^},���f,�V�Y�z���&ƳŌRm3�Ums��Q��,;�bn����m+N
X�f8O���8ӌ�ͳ�!Ɗ�/�:�W�ג�w��<��P�jߖ+\ﵟX��U�l%�J��n �������7���G�[��~T�\(�&�N>�u��\��S��^�Iq�£4�_#6Ȉk�W� �=ڌ��ǒ��ya�h��>��B9"��J�PL��<�	 ��2[o���^M���GCn�ċ_5
	�ksRg~U-K��_\�W	�dȶX $�y\�&h����N���Y ��n�v;o�%ux\[G ��I�瓤��N,Z�m�� A��|{_��jC��ZG�^T
���D��e.�`q%��
���h'Tk�_�"?�0�rդ�=Bd��9�m�1|}�'9jU*d����8@.��qW����?�B�kGN���u1���Px�?ؔ��0YI�{)koan^`���o�e�3ۡwW��-�~��߀� ��AG&����V`��I�.8If@��I��<���s(�◣��X��]��a�����7���P�w?~�XK�j��t�����Ω�n��93W��6ǾQ�.�۵W	���.��-V�K�-9�00����"��s��x�C���]2>�[��ͼ��)I����Q#��-A�^]������
��J�Y��ۼ�Y1�٠x_��X�,BrUDU���!�p���k���i%�H$,��=��,n'	1+�������PQCp��I]]���W3@� a��>���0n�D��ʉ,1���-��qCj�wu�^X��5�^����,��~C.��7��ú�o�A`9�g����1�}�F�%���ˏ�tZv{�$�TUy��g��?Е��7�	��E���gy�v��'�տ7��_q�AI�G11��>�͙c5�4�5������)�u��l,�"�D������b�{	�]v����Y�;�y&��{d����^�	��{��j6��*��.'9kxɊ��
8Zơ��h�`S{�m{�;
�E;��Xx�4�F���>G�Ӣh��{?p������n�^�G׾�W̯�/���p�ll��Y��'�:� ���gT���,��e+iW����f�w43��|b8�^'��N|��9!X(����Ծ[��Ӎ��܏T�yC��Z}�`���R�Gw��x�q&'YD*9�d�̥����opc�{�����ٝA��ʭs�.z��Y�r�<U�\�럇�xxF��g��n���k���o'�L�b���`��y�Z#�P���E;R��Z����aP�c�W�B��Ph}�m��>�ڝ{�!��Ɔ����6������	�޽�򪫕onli|w�⏫~g�1�3,�#FW�L�{r��tnuAr�lXʏ�M���u#���3F��~f����f��`���7��K���;�ߚ]���C����O+�z������� �8u�xc���Uc��R	�l���hW]���l��;��j_�I;<��a���I�`ʠ-�y����pں�%�q��ļ}��{�g�:;����9熪�Կ|1�A�&8_k�@�Bh\��P�V�:��{Mۯt2�iU��v�w���,��(��\Ri+��~v	�SG4�J��-`R��	�����]ն旝r��;Ocj�2W�ObG�z�Z�lh��.ɯ�P@2���׿学ԧ$M�����ۺ#s����C�F��I���NZ��6(h���6x���s�i]X��~�2Z�`U�+�,0y��5��m�l�|<�6���"N)U��H�?4����șc��u�������R�l���]�ź��ރ��б|���7��:vk��m��0�T�Q��y���&C���� (:���-K�j%�PW(�v���ۣ�jܝ�o�;�.�>	��L(�4z�x�[#�J&4�G�����ɜ��}���Pu���\��M�.�����e\K��
�Kxy��8�Ɉ]�!��q��RB�#��x�]�������s]A��'m@��`�� ����p���̿�ڭ}������(�(gk^PSg��7]~������5^e��h�(�.���JY�ݹY�zo��	q���y�s��-D� 2�R4�!K܄jz�|B�W����W>222vP"��r1ֽ�}u8��Y��Aj�������% 7�51���*毴�׶�U*�+�-_#B�eׯ#l4V4�4�_Q�s?ּ����j��g��s-����Y��=�p n�3� ��Y�I�Vz�%�Z�������^���|#A<ߩ)l�>�s��g)j�P�ܰ�����&��4?��?�r�/#S��>[�����
���5I�Z���t��������;�<r��w��#@yꎳ��w�I�K�}�T��k��>w�m7��'}�:� ���hXhYk1�כ-st�V�ش�K�XJ��ҭH��S�u��E�ZL-ϐ�=�5E�q�$�#��Kc�["|�Y�p��F+u���)���)�q]��w�x�̧J,��,>s[q�*�z�m����yI�j���r���s4詄��p�� 6*iߋ��V\R.�����0aj�	䥠�#S�Ma�(Ĥ�'���0u�h�i�i����u`1�5�ԍ9�s�.���v�C�t��v���g��t}Dd]?�T�w��]��{��@u����ZJ��}ȶ�<�Y/S��0���@[�!2�˧�7�<=��"���1�P,�%f�rHL�.���'囗�>���q��u�O$RPV��c�T����t/eQ��"�Ъ�Ҕ��ɂ�_	ǩz��1+w��,(R��L�G��,�Q��7�2���)�Mv��� ��!�'����w��O�Џ#�b�(t�r_<~��s���3Z�j���z�M�8�ֲ����.?
>�nSԫ�ok�ds	I�{���s�8���WM}���q�L�r��*�G�ƀ�"N�w����WN�M�F�JP5V��V�̃s�v�^^$�aʒ�˓�p��@�0�QL/�,�������ː�h"�[Zm��hN�ۭ7
w�{���i���թ��	�O�!�_2Վ�y����B^Z����[LٯI���W�(�]?J�ɕ�^g�v�EG�v��i>sC��[�R�Wr0Vs�ʞQD�*a�0�ı.f�a�UB����\�A(B�m�вݠ��b��|h��q��s	]QJ��HΩ�e�t���t!<�����f���`CO!��,9���oH��>�-;�[��
�eEٚ��3��5�ب��Tux��k����?`"�ݨe�.����Mb1�L#j"B��7�+?�����q2���My�w� 0����/<�4;u��>;�d�a߬x���Q>���걞fY���������J�)#ݣ�A�x�'��0�a�t�V���G����'n�����w�x�q
�ە��d#O������ߝ�m��<�"�8/�_�@��u�x��],D�����coF�=�����Le�"+^�?oD���m}C�z�W�1�K���!�@Ϻ+6l+����P(���I`?���K�ͬ��u���,q����1o��]��' ����@��3��%�U~!��B����\{`0
BW8��[o8���QmQww����a|�;PfZ�W��8�@A1������h $<���DC��<+2}���kh�N�<5����4
��d�P���H�T�]�Zq����C k�J�� ����f9��z���w�JU�t��-�~ �ӕ		�z�5(&�K�[����BP޴C�#9�L2�z�xx��BQ�{�Hg�X��� ޢ��8O��7V�d/����:���Q`g�`^�����=��A#�T��0���mՃ�!]�'b'}���U]�fީIO�s���Q�KRc����s2�U�Aʯ��}�'"��<���"#���z_o��WEb��C3�pť��M���J,)��P��XK;��Sl3f�6�J�PH+p�<�cp����{�Y�7$�u4@=ojյ��h�҂�N9!�k����ݡqzӕ�T�]�-��3��튲�T�3-j�����a�,�K�������t������KG6���X�� k���p�b6ƀ�sR�ˬ���z�V]��K��6#��ф���x�M�Y�����
�3m������Y��=�TH]���y�څ�d�2=�4�ғ��6�fD�~hWⓉ+�%�(k'�4^m�%M��D6�\a���0��	d�N�J��k͑$g�X5
�ݞ=���-�T>t��ǩ�����4��_-@�ɇ��
�Ƌ<��6� �n����G��G�B�PP���W�ܞw[�S<����q<+<5FX�H�����E|w���9��ef��!>������-Zޗǋ��n���GZ�5_�� �Ʀy��:�!�����C>�X^	�;Zx�%u	pB@��D�yi6�X.ő� 1�s�Pr~������0�?�v��-�p�c?��=����^4"#�`�0�<ã+�:����k��_���])�qb�5�O�䕆��0����hj�{iT
�{�n�1�o�;��G~�`���C���p�~����P-v|��jQ�҃�DM���@�=�1F�~�q����fw�Zw�i�[z��5)]�7��y��3N��)��E���#ꭣ����q@:�� "�ҍ�tJ��tץ�A�����N�KHww�����~�\ֺ뜽��<�̳g>��!zz8.RZFw
ؚ���=l�S�=~�ؤ���ViU�o�(��[����Z�g���65���ھ�?c����֨i�$;���K�����WDxڷ�]`�<W!i��[��o�o��9S�q;�P�0)�Wz�#��j�#���YA��$a��0b���M�{E"6���&K��Y��t/��1W�tɗ�FbU%�����)�C�,u`���
=>������o�)F��cKz�ڰ�ȶ��d�	�g \��� _�]�n��X:��J�����_�)+tc����S�ɪ����Ah�x���dg���]`��R�1�� �B�G�F�������T��0�w/U��g�|p���,
��b������`� 益��\��7S5TK��QȂ$�>����D�Z�ϻ�Q�a	>�ɳ���E�i�}��'����%fWa��,{����`w�(kDv���	�K7�Ph���޽���A�^�%��,3���6UA��Q����^p��ڞ����L�iJ�j���Ep�@~�A�%q�~�Ulls�7��u��t�T�(^���@x�Ӏ�3�:�nz��`�o�@���٩�����P�(�NM��3�\���L UpvfE�A�i�5����sVK�@��e����0��;�I���g���=We9�U ���8S�Y	��X�/5�'�V_q�p�v�L�|Z5:��s�¾;0��8x��~K�����y���Y�����]���V������?u�\����@���������6Q��w>R��\�x��\O��J�iڻz��k[���0����E��?E����W7�T�2K�F��cN"Y�C�%�\2�Y/�^����Q��UH��1s��i�?�~-z��E�{���w��*`�l�W�_����.7Kl��B��J=Ijj����|���Ǝ�ǖ�������ɘJ��@�U���N�p���d�ˉu
z-F)d�v�{��c���F?U"5�c�wZ��1~^nL��#B����(�V�T��:bOp�fdg�-�[� �0>Y��ip�l�������
���$���}P~M���*��d>��C� ��K9Vi$��\kS��6c��q�A{���&��ǜ��<�e6�މ�ы.�ĥwgV�t銲��GaFҭ��=$�i-	�+�+1��p��R�>ެ�oɟ:�8מ���F����l~t��?�}7I�����kv��p����x�4��a�|�c���{FOI��h�����%,��S�gKGr|�x�m�me���W����h��?=+��j�t�&�{f�}��B���0Qz���'*�EuI8i�f
C����0���%���j���L�>lĈ+��@�xS�'�
&|;���5Cy�9�+:>.�2z���w�=Na	�K��;PDv�9��_�E��z'������E�O!����.y)�`��B�~� R����E��ܠ���D�\�3�e��}a
l}�$��C��f �]�R����=�����ԯF0cv3R	�_&7u�]���Ven��Wp�찒�<�W��:stKR՜���C}Z��$��Wz����v?��E���_��?u�}�|9Ϛ�!��O�׶��Mnz=E�;u6���ֱ�;컨ٳB )3�S1���|�Z��ˣc8K�2i�e�k�o�&�'����ir��oS�}�lF���`�ɀ�a�2w�`�}�VR������jة�w�W�m.��a�>�o�R �;;>!�d��+Y�_$""�����F��_�P�x���P�L�-���kQQQ�k����c6²b���jf� �V�/��ퟛ}8z�j;OF��b�7�cX����������%�1���;���ВXO�A�1�mZ�������׼�1b�6�}�M�|��9��6�I��0`�>��W�BYNm�p���HE��l����i댒�Q�O��*"i�Ob��|��k�����������Pii��ь�
l��e|f��	�J�Ji
7"���|��(~(����UC����܈��������E�����e`��
��^Pцr��	�{�q| mp���m)����a>�U�t�~ӱ)�
|7VPLd���K�E�������CV�(.$w���>�U�@s��H)e���$�a*;$���N�	�%��^
�rh)Ƒ�g(�����@�����z��i?��ؘqѡ���1����֙3F_+�n�lti���]�=DCMm��I< v0}�R)�\{|���?5�4�C�qؒ.���'S<��ܘJ�N�]���cE���2F�]�s<���^W��H
FTL�\k�	���,�|��+��$� K���mi1B�ii~>�Pr�뺂�$pf��G6���A�iȬ�FJ
�T+��`�n��vzMU&")���/�\���L��#�Jd���o���<�ҷ;�!y�<D"ya�'��T�qC�&����C�bF3�����&+����S�G���~�!�/�h�H�,�$����Z��|�kz_����iX;��b��&�ƪ'E�=��x�4��eV	U.��mQ��̗�u3��K����=9m��ߔ1�Z�p
�4(��f�Y[s��`�X�h��-/\�Ea�jq�� ���4�]`�S�k�M�?f�Y#Ѵ���i<g=��%1z��|,>Vk��X�P�>�@��hAj� ���b�G�U�������ƒ�9��ׯW��.��γ�w�������Ҫ��hR���P�\BBB�����o��&&Vu����`X H���z[�]���^���}5j^��8����|��U����M�ý���8&���5�Cw�Y�8#F?7I�7.�1DXIQښn��Gy�4�]���~ge�S둌����(��"����U?��b�����9�4��&j!��nu�[V}4	�$J���_H�H́���es��8�l��<�17	TI���[[[�}PN�䢟A,�MU �K��$>��D�׳���)@��~��d��R��VY��*S��͠��2ER��Ҽ����9��\�D�u��n�̎�?A5�k+%+�/G_���K���a�/�L�c���⠳R���GU�;�ýB9I� HUW�����<'� @F�����*�������Px¥�ځ:�՗wW�<3�A'k�o3���c�̜���ol.pjFC�oC?GT�.��L��z���^�=86\�a�W�{uE&"n�X#�8��9�H߄q�5�=F��ڳ�~���]�a]�E���z����)$	��X���7P�����g6Rw(�x�\,�av���xR]�� �o��
D� ����+@�*�H�3�_��kp�˜x]�G��RӬQ��s�p�hr�{UC����AU��~��d�wKk�����m�K2��s;�o�>��|�#��6|�nUg�iv���@�'C�<���Gg���d��j�n���]M*��iϼ�apĮ��f��}�t�
Q�ZA%��b#������}��0��׹�kc��>�V]x����*�������ժ�m�ݖ^S[�K����丫� ڲ!k+8=|��*�Ę�:�9��3����H1e��$C��8�8�q��f����?��*F��پ/������ջ~��]C�����c��S}���2\Ҡ"�bSF3�5���DE���>�-��	;n4�ݭa�eV��^�n��5�V%D�9��� r�|�M��Zfw�Y�N��']�:)�+���y�Ar1���;I���E���9+ƛ��(�z�
����!a��e����n���=u���cg���jwd�ò�_�n7YЃms�{PG��G�qs��Gr�ˎW�<�ʏ�����£*�_r��Լ�ڻ���2 ��Q��Cp���!�&$H�g*���
9jW!���Լ�b��+Y�
zuU.F Lk:�<4���&����e�6��g�	�}^O�j��`*)Cc��.YQo�����2����}�OoKqh)�����۸n(�;�ջ@�~v�\gE6����Z�\��us� �����q|D[���?��Y��o��r��<ρ:��fqG����e,� �	LH�q�g��-B$����k�o�<J4:ƨ̡�nʴ5�b�!�m��ݝ,�}���e+ßBY�1�\T>)	�n�5bj�;!r�/-���t��:�^�|�����e
,g)k�{2ތ !q%�L`ECA�	y�#-�Ul��®M��̈E�V�x��
�{��u���\��jW�4ݤ4��l,>a	b�DP�j�?��v`��i�����a�^L%�;	b���Q�ӚX:��Z� �D��/�Ò�Ҷ��99��U�L���D�eK��g��܆�!��!Pk1�mX<���p7�k%jj\\0Ĳ��
�������������Y��*)Q�;�\�� ��旰�*�9�q� v}̢o��y�6l�Xv����jF������]g,��U~��V��bcq��9�iz��]�]�Tn��N�wȼ�
M�R�i�9V�s�dΦ�\/ߗ�u6��허���+��Vt� �,��%��вM�]⎻���G�[�ʹe�Iܖ`r�+�A�
?��'��[��y�<�]�B�[�ފmD�IX�-o�-����~�4���2fFO�3NOWf�5�lU/�N-*����?/�Ő��A,$H�Qp7��10���I�c�}�GQ=�Pʬ����][W�z��!��PM.������ʙXx������9ˌ���Ē�V�!妖h�nY;}��>:�â�;����d����fd���QӤgͳO��Y&GlY�-'�C��$���7�8\6�N��<WB���݀)���&&�`�l�.�D��Qf�Ƣ��OWB�d�o0*��3k�K��A:��`8Q��n��^ ǭ�� x���O%a+uZ[�*�z1.#�]{/"@�G�hĀog��n���G�OJ�������R�>F����A:_C���<o�"y��5D��5N��7M�0����c �po+��8d�����,e��X��A�yϩn�@"U��F�� ������:_���z�������<�De')����f�=�>֬�e��W�#��#i��.��Q�ߤ�Q�tϚ�l�O���T*̏L��\S�ԉ�~\�Fh;-	Iօ�c�qp��G<Ǩ����"�g��52�蝖nF��w.>�li��U�
��������9��wn�	zm\?��H������ߜ�`����O�m���|^3-��L��Fh����{��'�(6D�r��� T���s��4'��<{v��q��)�6_�e��<<_�pE�Z��7xm�z�[�m/Zq��\i�/�Z���:��ۚ���g߽�$f����F�4�1��Wթ�'��w�?��0���r�/�ǡ�b
/���ql����=�%X�ݐ����j ��|Ps�Je�#��;�Ɛ9�`2���R[�)�tm;Qo����~]�4�K�K��eA�E��F�-_���3�{ktؓ�����/W<���	g������an�De� a�n�fJ�v:����3�,�	�
��;�e�����~\p��K�a1�cyL1$& 7E��ވ��b�@/"��&Wg�D*�����t�k�}{E|]��*ŷ,r�l�\W�H��Yq��s����q#N<<<�s�~�7g[`9��tcp���B�b���氤�9ܖ/��	�TH���a+W��*��I,�a�Y���텣�KY�֣~��"���&�9��(h��#W�R�+�.��Q^c�b�H1�8��tAf2!%L���9���R���"�Y�;��+2�r�4Y<0�Wʜ�߷xP	�h����T8�����D��U���>�^��<�
>�� FTe9���*\����7	��%~���`�A��jwߨ皵gQ�tP����m��fq�,�Z��xA5X��UX���[���+�����c��>�90R�,��,�D<��u9&���ѣ!ٜ�H{Y���A�����>yzt����p��^� �c�J��� W���+�?���Y�1}���s��Ou*�����CG�y��y(\����[q����
���⦛�,��)�Ex�����I�F����x�q+Nu*L�jX	��4.��ٱ�Q��U`k_~��{��u �J�,,]��p ������ϯ|q����>�y)�k�����m�s�"ˤ}M�"�,&�;�
��,%($��y��g��,�?[NMz��3OM�8kE*�a�NI�Q'I��8�P���אE��
�&�tm��(L�
&Bg쯹�V���		6z�#��T���ޯ�")�_p����	%Ѩ��u��N�����|8��h�ݛ+��*aN�j�/wB���5Н"�r��ؤA*�O$��)�`����(` ���
*@6���}ç��y3ב�}��%is2���Y���s�����5m��9��F ���᲻�u�xj���o�EHct0���!�
�U�ڌ�
e�NL�P�r���D��=J,Q1ҳ�2P3���XA� �/�03��֗�E��!$e�9��[?w�p�0w�
 �z(Id3�� �uX_������w���3�M�nG*�d
{�Lu%ŷ�%ă�|��!��:-&�R6�/������5����LÍDF$�߬�d��k��N8���\a2��HW�m��H1��㕮_Q��j|{)��KPC�f��k6�Z'k�`�7Z�Æ-��P,�݂���#�t��$!��G˔ �_�[qo<���I�_�΀�h����;fl��Qi�&F`�PW_�ih֘�+��]����Aٽ��2ϒ#�$�F�P4�w�g\�R7�z�K[�)�8����Fv�"6Y�o&W�s-Q�l$�
��-����>o�GT��ſ���趤��L����u�N�%�S�u�~��]���N��L �V?[��:��R��s�$R����'�2�y���)�d2Э��#�'����`�N����E�*x� J����6�aར�U�s$���|8a��G
o�G3��nFS+4P�"�(Y.���Ė�C|�u��vGW*�rGS�C�ً���F�v5NY�=����t�=��
,f�R��� ���Nxv27`+�y��"��o�P�
���HǤz&�f!]'S��>ajv�$�4/��#�	,�y��[���hVP�7
>�iV�q<]�R'0e��K�$��f���w��_��FV��x��r�(Lj%����!E�/?=,�9PhY�S����;0P��������1s�=�Lv�T2�o^��h�I>p��ٲ���7��-��
Lm�h��S,�9��=��s�Iɖv�� ���jͪ��M�:s���*�B6�'y��W��o�K���p�
���$�`\i�ؗ�����A���t�>���$�v�m���������*�y?�A0��	�do	�J�>�|[���� ����}!�{���&��'�z;�$*��~֋-��hn���&��y�����>8ѻMC@� n����� ��ӁLL冞7�y���@J��3�T�ߔy��O�S��
Y���Ʈ05�J�ɀ�n�:e��qH�����:w�zp��G��w~�҄����|Gf��] {�<�U�7�45	,Fӣ��#N���2���������"g�R�ru��n��E6��m 5Q��%;h�9n,6H��fƩ�j�ۑ��v�Uճ�#�v�+�Hݓ`$�	�Ǚ7P।���vw\�Xr�-�)�=59���Ȼ9�Id�	����Z�˺�����^ as �nMIkkSrVx�x��(�y}QFo�j<ﶽA&���Ju�$S�����7����۰��A��2�/��pw_S�@=Mk^���5���2eT�}��@����:,��,�zc}��	�f�f�T/ܿ^a���r4I��|s��T��?]8~��el��S���p\hp���;�r��߰*�r6F��,e��7-�v�ڤ~�ԃ�����2�WݴZ���\_�l�/�p��-m�a��)�5�7��ؼ����F��w��j�d�U=�*��Ab���;��Z�	b�ύxÜ�~<B"�sRs_
�T�����}пhjj��3�?W^ic1��wu�^��&��S�����O���ah��ە�:��U;h�x����nFnU�e������߾�$�|��4	#���!��M.�����i���Z%�
��>O\�D޸#K�&3��t�%P���k�=M�Q�����Zѱ_܄�Bg�CC}��|��|�T ���,�F�������X��)Yn��f���`j��a���v�_غ�� lJ�� �WG_�,���� ���Y��3�TDn�t	6|ߙ�l�mْeҶ��x��G���WU/���<Q���������2@F�(��y���r�ߢ�Ҏ˳�o(4�g��!����¢%]�Ȱ�1^��1��⧟�p��)m@]�����ѵNlQ�����\=X� �8ؒ ���<R=T;��"�ˬĘHXM����5R�3��¡��@Y�i�NM޳�SZ����D��j��S��I���(��1<��C��[��v�+��"tL���
�u���F�(�m̻_z�Qc�a�^m�L.ΰԶN�~u/��,^bĂ*�4Ψ��oI�RG,�����{���Hr�dhr��u'$��p)+4�P�%��jz��9�&�S�!���XA�Ʃ��D�|��}E(#�{*e�}B�^�e)wE��ƺ9DS����)-:�/��6Q(+&��i�'"ۍ	/��
�F6
Q ̟M�a���C'T�F,�q�Igp����~�S�[��M�@x��{~�Ł�mrs��J@�g#h�CW8�O{��j��&��r��*�����ޢCó�/߀Y�{ȼd�J�qc�Oc���w�4��u*J�����n�a��!�A~�z�Qt}"Yf��;Q�PD���j��c�	��p�:z�vW��)��J�|a�=r����,���tm�E��?X�ykO��*u0ʡ�F^�<2�}bAw`�#�E�Y;5����сQ���R��g�9�}{�U4`��$��������Kv�|�:�s�$s�Χ�ۤ��Y�֣��:�ڰ+�_��gX�Q� ��T�J���I}D��᯶�9���H\�ѵƄ[�N�^+@�V3�&���ƙ���*ճܫT�f8� V�i���Ov�Z�z�t9�B�`����.LW�>'�
Ŧ|N�M��W�Ķ��>�4~ɝ�=@>��Fi'*$���c���:�w�p�%�7&j��8�(Oh���/�:18�!z�:��a<��0>�;�a�#!�WU��P�?2������r�i]���n��`��K���"������>�<5q���#x��L��f�y��A(�=���"�������P0�	��\\\�}�ƚ�p7��$�)2�r�[Ը���~a;M���B�� 9����S-��Wu�ce�s;�O��o0���kM���/l��Z��G�_Ù�K0����X̥�i��[H0��Cg�H�AN�q۷U�n\)0@ ΄�7řs��k��өw�6�9�c ���lpն�`�_�W�b�G��	��;����
�*ݑ�����Y��?'�a��Q��-��J����	?vLC+�-�_mb;a����JD|������S�a����c����ή��M{���������oiM~�H�%���"Q�Q�Y�(s��.�G�G>�)��ڶ9"�4;�>FCX�i]���2[��A�5�@�~����v�2z�2��Zc \�	+)�E�����C��of��A�b��f��)c%@��S�1+הoy̶�RrYe�������V��5����{PO&���Ʃ�E�C x�W�G-T핧��f��c�� 6z�qb��9IG��yR[�Gx&�@���<ׯ쬬�.��/)�����3�2C���������, �����	)�������\�Ww��>��Ԋ$�u��Fc���P��������u�V.�e7.��.�-����u-c�42��H��k���X�:�;� @g$R\����L�����ӭ��C����W�a��N�j^�^!Qv�V8�G���L��e�����m�x9��9��Ф�0뇆�d�P�ƈ�F��8��!V)__apѯ��)����mo�W"߸#4�(�>���]�f�����ݚZ����Y>E�
/��xӇo�� ��y���2��\�^����_�8��	���C���qK�%j�*0��P�U^f�`��n��5z��4�_}�snఞd�����乆ŢW�)�q�c���AN���33`C�X��/=.]t���.����y�����f?��LB��x�c#ݧ�z�#��������R?;�N4���Y��'��EO���%�+\wt~8���JD��~ʢRw�4F#9U��C�Vֿ=�����s����5،߆Vz0P���R1T�n1!v�6Xʈ����}فkL[�bCE �ρZ��Fvph��`����1���9(`UJ��"��W
8b�:o}���%����W6��?�H�`f�b)	&t�ϟ����P�j�&,�Y	|���+q��S*zp�kʟ��6G�Z	fA��y���+�4F	f��ψϚ+�j��|���Ls��IV,Sk��e�͎S�ڠ��s+ͣ�v��ب������Z���2�h�-- 惫dV���#�fdv�b��X��y��i�VW�J�ѯ^��c�N�p�c�2���ee4�լz(^�va�D��ED�i��Ӵt�/B�:]{V���y�eo��z8T�-�L��=G��B�@>��s3�>�љ���-�[�7�(^zv��G�x��h��,:�pg�Ý��/7�Fo�;l<�@��B��E��tw� ��Q`�7�~��l�4�4 8y:�i����2C[��V.Wٚˋǣ���o�!�� C���=6�u��#��ы������֒�)�J�]��ޘf\��"F�Q.�v�.w�2w�:�9�:[yMg5O��k�- ������L�.��B'�Ee�h �2ddc�	F�g��������z1�Ü�]��5N:����`c$��"	Wp2�k�}&�I�.&칺���6U���T�w�"�w�`y�AI:�t�[y��� H��ҽ��m�=���e�Ne�v̿����j��)�,�B6�(��&i�5���$�k̦g}�)�>�Z�%��������.��!�'�Z۹�$#?��s��do��'0p�%���;��c">EfJHs��̏�>LYJ�~�d�h�ńjIA�s���� ʬ��\�*l��3�_�K�mc�<ۤ��D��o?g�cr)m�[�!XM��\2�	d�DH�jR?'�
'i4�=`q�Ͷ�
�s�}�4��`D|��x�����}���'z�H�(���C /HĽz�q��g�¬w�~ܧh�N�k ���]��
O1�`�Ʀ����IզQ�L�c�=��X��'�{��v8�O@8��S�5�\j��Lį����!_�������'+�C[�Ow��a�'yu���Rqu���u�4D�Y� � �c
� ������1c�L��6��u���sjk	떼�K�/߃�j�Zn����|eq^�;i08bƀm��#TUT�\�����*�O�\�'I�	ͺ����c��1��r!0,���!�N���� � mD�����|�����M�g������E�������`S��v�Ě�x����E�8X�)8��łEٹU.����� c(w�RۇXYY�M�譕* �JIS����XB��k4�T'd8h��`���o~�?̸��CJ��W�_Z(E�E	���Xc���e޺yI���r�B*�?G�J���^�t�*יY�R��Z�F�V=���r�d/j-p�]��{\S���1�1�+�xNo�Mw*�"#��.H��C\\��>4T%MR��YF���R�s�Yp�:��VU�Ȓp[dVT�i�t0�56C��m�
������������y�ݻ�Vm��FmI�.ڷr~<3��d��ъ�X���B^|w/����#~��]6�U���>��qܗ��KZx2��@����c�jw���޵���{�YX̝��%b��x�i�p1?�-��^��3�Q_*��)������CJ��\.���`�w�@
������Z/�An"z���qhA�|�7Yk<�Y���q�k�|�S�ԔyUl�J��l ��M�ܲ~�ᯡ�~ĕ�����_ ��
��p @������x�Wǉ`�L ��y����(cɣ�&�+kmބݰE�8D�@ԀLƾ�o<H���pꇅ�b����$�M4����|�ڛ��3F_�I�YY�{�%�66��Η���s���opr�~�]���1�<���#�� ;"Xx������H�R�:�����F$��c�/���..z_�D���`펃(7\���VWCEL*3B88$��!~�_&� ��_�c�� ���!܄�KRYY]�g?X�����)u�p�/sZ���a�������9_E$��PL$di�K�`��é�R��U�\Cq� ���^��śƯ�5��{�F$|u�5Ҍ�NL����ӝ�:愎�%�I�DYݔ_��p�<�lŌY�������\�u;�`
ͥ��(۷��&�|�)��]f�{c9�{oBB�Z���f�:��_�٤~}�����d�F��;[a�t��
���P���r� ��	�-�9�?����=c�W:��(L͗n���մ�3�\���tG���ś`3�E,~VL �'�;gg���d<żԵv�JT4���+��u����R�>���!��#_���;;��&0���5a�����\p$���̀����<`�9�^�D��s��z�:A=��,�e�������%64�V�)S��|/�Q��x�b��`���9��5�Yi'\m�-:���U������1��］n�	l�	Zb��&�du��������dfE5��+x�Ӆ[�H�g��������(��La�u�:��=�噧����4ع�׻�����C(
6�O#Y�����bu����HD1���>=�Y���`-�������!~S����:�S�%�@��&��2E"6��Y1���5�5�ru����v$z�u7�[�rMCAa�-��2��R[Gmt튞+�z��4q��	�E$q�HM�L�O���Z���#�����T�T�~��]��;����`"x$��z��1�nُp@��ݘ��%��444���9����F��� �ɮ!����n��8���0�Uɰ�]��������h��}������U!����K6��~k�9����S�2B��e��P��£�����:U<��N������Jy�����|��-"��F*�|��"YΊ�t!���t�������*M>X�\�i�g��"�����/ɴFs����0�9��n�'+a���L	��v�t������j���񜷝���s����{6v6��oz��L0wW�^u[����S>��c��h��Y�s�����~P��Yu����9%���6�Y�l�<�g�膳.F)��i-j�Z1��eyL� ���@M*Y� �~:S丠�Q%����]
�J�R�Cӧ�0�N�l����ޡW�����E�CBB��'��g#BG�Tu_���W)��ފ���%i��
/V�^�ޅiW8οw�&'}h�"ߖ��Н�2��?n��GC�y��Jl��*�`W���v��#��ga� �C=��ټ�/H]��P����|�����^���B�W�g/�D�G}Ԩ�H^͊��L`Xg˹@��T����z)� r00��a��J|��%i�2�lx�j��E`�^{l1��}����ډ1�ܜ����YS>]�������d�z�Cp̥ d�RD;	6�a`eE��>��xF4��]=�$Ur �z���v���#��H �Y	j����^�?%��)����;����?L�K�Z�5��Ϯ��d��	����G��� i���$����WR�	:�3cp%b!}K簅��!2�g�Æ�/y�_�P��8R!?'O���F�k�����}�h�&n�������*Ҡ"���`��PJ�|y�E������ŝ="BB�'�]|%�# ���3����o���-��D�\���a��/�)�[)�كM0>hu�O_*V�ǻ�Jt�����_m!�f�Q�u���:J��NR�����\�1K��	Y���Zz�A��:��9޿`�Ͷ;� V�U5�Q�U���¤!��ώL&)�]�6��=}�X'��=m��qpWtr��4Nk=+�0�N�C+�iŬ3��AX�3��ҹ��og*DQ�h�;�=�������C C�A-�`4��*>'ܿ�p#�;�$	�M����+b��lJP#�N�������sC[�\�xv5�([K^f��%����9�Yx�F��븂_���܇Wh^T,������ld��`�3^�,%,��sٰa�����UI��pX������S���t,����H��B�H˽/���P���) ��N!���LW��0���O����i��Ɯ�>L,w�-�ʈ�p?�<EQr$nG���{ɘ�;��^mŮQ
(�X/�����+' ���M��Q�������لs�>��憎���tn��:k]�4��/���>�YEƮWI�^C�\�R��Jv$[�4�A��ݥ	�=�J��R��S���ڷ�t9$^9����c����B��G[CF3� v�T��l(.ao}4��P�G)�����J�8�u�]�����F��,�aL�<��>�{@yy-0�:%�@�P<�B������agAb�V��$*����C&�9q�YrY2W�Ϛ?^y�s����x�(@�ܑ�]���?r2��B̥3�`WOs�goD5���bs��<&�>��R�pP�2Pe�G����pG�純���.=�_kZ�^�D�@/S�Ⱦ���g�{��o��s��B���ÒBh�������֒Ȗ���@̂_:}�: -�$�A)�o�VE/E'`��Di(T��2��ϯw`KhUmm*O�������ꛜU�D�g�ӈ�t3�(<�P��r���+�D �y��b�Z �7�z2�K�+l4�@���i�+���%�+Z'��EG�f���P��o�h =��&��Y�'�ޓ��$�q��fv���2��,�	�39�ً˨�
���ٚ=�,:{a���������:�����
x9 =u�+����D�"�X"e������[ߩ���t�����n�+�p:x�wA�dy��ј��e[S�M"���8>s�Iz�&���ύq�ɳ�2�3�!�g����[+	�yN�+���xů�#�������ƻ[�(�{�^�.$��/^�_�xE��pN�f�U����+��{�z�)�M���u���S��V<�*|I
;������H���'hmO�=�r�����$�޷�ς��qO�t��J{Ӎg?x�����9����s1��0�LT}��R���~7ˍ�~��������	N��8x�2=N����<�<�p>k�)�S(-!q9#�<�׺��m�hB�c���g��*Kt�,�?��ͳ�E�Me�뤧H�M�3,�hͭ�=ؘ�,(�}�[ׄ�ܪdD���oKן��r
D��5��
5=H��Q�ӋN�[�d��N��@�����d�y�ls1v�����|��b��ڢ>�
s7�q�|�;�3Ɠ��'��i-5�$>��j����=���$t�_���l���Nͥ���b��}�1f��4/�*	��ċ��\=7_*�GXf8�bd�~9��Do����^��a�yL�����d�'�MH6�j��H;8g U&���BZ������L�O�D�zZE��{������q�G��$R�2u���Z\��Ŧ* �"!$)9ހ--8�|�z��({��b9����Ho���̍G�箳�
��)��~��fs��_[��@�t%ɷv�рQ)����	��h$WJ<+=K�C_�x�0[�j�%��<\�<�z�?�-Rͺ��]R��
�?���]��*�2�繽���m��*�)2z����+8���`=N���3�!�*�A�1l��\��8)|2ff�pвяK%u[���E�R��g���%nˡN�e6��勌��X���ݕ�8%JP�!s�|k��}���78��Y�=f�4>CI�	J��&�7э�J��P��<������4�D�Nn^5�Ҁ$�fK����"A�{�lM�/H��Ӟ�.����;;�`�*�QSX�8|��W���1�%0Yzrj�`�����"�B"�fS蟃�5�J��!r���53"}�4FV.M˅�%�`�fJ	�L1zP'�V�Sa��wVdUy.���7�0�'�Qؔo�\�bM�i'_��we���8��;two�T{�����5:�z\^=�#��=�Qs�S떔��
]#�>U~"��o��P?�]��Ib=�������m�X6���pa~�c[`#��h�&�t4_����ؐ�#)>�C/>�,r�?��/�	24Kw��� �0�d��Ƞ�
��.�&�^ҕ�PY�(�����Md�%��%y�eލ3FM#9{������ub�ux�%�!����ӹ�0��_�T������A������ظQ�Ŝfm��jv?^���f�,�^X��I,~ej��:��f]0�l�����>��-�}螝�ǒ��V�f����`e����E�Z��ʢ�k�#���b��F?q����@x��j���Wc��,]�ćüۼ�>�d���`IWt5�Ftn�y2%���[0�_�}g��h�-r��V�F�8�e){2H����*��.j�9z؂~�K�̞�����rd]�oo�"��qNξ=ݑ��I�v��~c��p���?��I)��πW��������:1�����A��5�A����������yoC��UTk�".��x�X�uf>�;#[F�k�g�v �ԕ7�?���ɰ$��t�EJ�����R�R�0B�� D	�1�Fb��ݽь�{������������u]��,r�c�-to�r`�-�+��%K��������׆nC��[ ��3JKKw�^0�e�>8	����tIC��U.iI�)0w�W�y%as����L�#O�,�,��H)6��R�sϫR*�G��;Wcuԅ��u/,�E�ȴ����Y&�;}���I��_w
w��g}u{/t�c�I�Ȁ�(���>&|`x:h�.f��Y�~w����?"l�v�qMj���.�s���R=.��p��U� �Ŝ�r*�(����;�Hoz�9�O��z_FkT�*Ro4�ғ���"�����P%��D{�l�E�A��E��" =i(o��&�ZN<`}Z���Ģ�&�����\�L遆&œ�<GE%W�e����%V�t׷o��t�/	�N�H~z�*�=�c�;��#������MлW�5{��7�����4��d�"g�O��� �3�*�t�h�+����Xzϖ����1���37�U?Z!7���.Z\H�{x�-�d����Qū��/`0���isoo�L��&��aMq�E�`uN‏����Մ��H�5ت�ŹʞF�l�h���[	�NC�(�d��P�%�~��o�$��ݽ�z���6������}��ʸ�n�\Oi�1U�5��/D���Q}X�B��2d2�E�΅��0+��.����j�������ܥ���v���q����X�����Ǜ|$qM- �'q܇�s�ta�u�'2p�Wz#7�Le��RUh���]Y)�(D��v���c[.aI��w���}f��`�7�z3p	����0�g�oD�&�0?��[J*BI
��IL�Tz5y�qC.s�颤�_�R�y��.��%��W�am�Gv��ҵ���~c��X�&G���+�{Q���c���ez8�ˎ�^[��+���1�!ɪ��h����Î� j�G�g��su�n74x���ޭ�!����l��/3fbǇ���J�tc�#-����t{ܟU�#���ٿ$e�\#���mk����rǙgEz��qD��;�OOBW�쭣7X+��dUg9��f&%�SX_�A�`���8 ;�)K���ȁ�<Wuou}O��H�z�.
5�a;o�̳�����BĦ5^S&K��nv$��h\��3�2.�NZ띒�("d��U�_/Y�����8ռ=���8�,�L�kE��&������N����t��kGG��P�W�D<o<��s�Vrk�[1^{���w~���>'�]����C�벨5�o#+��Sb�]�8�MCzl��	��i�V�k�����'+���K������9��3������WP|�&��/�땝gr]���`�[;�$;gfԸ�_���`�lR��=�FG����d�5�|9��֑ˇ� �ѹL�(�����#^k�߀�L��|$se"A0�$��=c\C~�uuą��1��ٙS�Z�/�M����rs"?�K�h���%��I��s�I�S�%��B��<j��N�AIV�E�[z�����Z�������"�;B�	dweq�|w�D��9پ�ЋYX��ż%]�۬x�y)���ꢤƷJL7w��`��{Į��`�� �,�+Y4��YY�gZ�@�T��Zaa!n��~��O����T-����|xX�7���=b�;�ڥ�h�`#�Z*�m��(��`�����N���17p�m!��Q)�q�g� R�㯏,£�ƀ�φ.�!8N0U��	���^(�m��\'�?�P���]c�h�����?\�|B����	g��ͭ�Ƨ��G��b�Ճ�y�Mw�O���y=��0"N�̫��Hk=�~]ҩ������I�;t,�cҫ�M���JiB&��H;�̕����`�a���"y�ƣg#g�k��1}�

�W�7�;ӎ��Y�͕�~0 �;��Yd��&⻯p�R��5�pq0Ѕ#^			��IW���L%��{E��z}B�.<B���cPd"C����������sq�@�9� �?T淰��b����Vt�+>K i��ȧT^���?�*+�/s�ژ��L�e)Yb9�苣�aH���ȣ��|��Pa��s��颣�J�;:v�$���t�DDg0���j;z�L�p͵��p��[���33��
@��Ą^��A�&u�������I�<ݻ����{x�g���I5�B��e��$��Ջ�<�Q���6]iR��`NH��$�J�x�����$����xjtַW��d����|���g��*ǂ4H�5E�Ip�k���ja+��&�k�G��W��`�¿�9��c�ůCD�_@��)�@���m�/ӟ�ݙA�VW�����>fD�����	<��.i퇹-ގ�P�`0X��Lq��K�g�?��R�Q��ǝK����lY�+�R{5v�aL���GHr^>7iP��L)Gb	 .�C�1��="]���:(涓o�>�I~GT���HҶb<�"J����o�:吨�����eP4$*��D��$8��R�<R@^iy�55t8��྅����$	ô7���Y���5�޼y��+nxb"�����p!΃323[��:�+�����M)�<�n�	��v\��R<���^��OK���h���j�:��Vt&��nI�b9���s�ŝ�נ�$�N�i�ެ�<��^����.�}�j:I˾^'N����z/�q0vM��y�(ztgG���$�3��n.;��2�~�vI3��	���C���ԗ%	�W����.�}o���#'�fz9�0Ш��-�ƥ��h[��;k�L���q(z2��8Z�����(u�!@ѵ�`�čj�ێ�6.?�50��b��,��uu�JD���<&��}�=��ZP���mm/z�i�����O�3N�H�`�L�݁�����	 4А���>�䥆�a�m9-P�M�+�oo�#���ԯ�)�m9b$Z��hgq���]�&)��܍g��y�O*���%s"�6�2u�a[ �a�.ۏ�e�Ɉ�������7!��s�Dh��N{��?1�[�YK��ޙ��$]dX'\�U��>�t����ר}���&tf�S�<�{�|Ձi4�L�����j9Qa�x���bp���YJ#��[�28;u��ݩ�� j����ׇ]��eŅoޜ�p͆m]c�N�'ai1I[ާRcK��� �^�����0V�L�{IZ>�q:jq]W�q�}�����N]��>�q�]
��fQ��M)ymM����.�CW��xYK�{k��^,��Y��K�}��`�����QʂH�D�����x�e	�����Prֻ�qI" S.)��>9.�Uۍe�����2�\��>p�P~\z?P4 ���t���� ��u#3�9��7�prb�G��AZ�_������H�?�?�4f��Ru�"��f��Y���￞���%$K/'���3�N3�/P�]�{�s���涤')�q��x	^��c����'}Ώ i�m�N.�,��@��A�Z�Ό35�m�[�]H�$G�r�X�0���TyE�����#1^��z$�~�ߣZT�٘�O�����G��ЯJ	0�@;�K��dK����#�&�Y�M�F��.j7n�_��P�PI�
O}{m��h<	�>�n<u����
zg�@C0}���Ks�(z����ZѪ�.&�߷�4�����3]��hd�h�k?��@�{_���ge���(�Q~��`�ԗ:s�e�C���@�
�6�_��J�i��񙮁4�������M�<�B��Q���#�p@�Їyܔ
 �Ē3Jb����H�ƞ%�5<<<��"���Pk��8J�^mRz��0"e?�J$ć��$�MEM��LD^��V�lv)�f3��V��fj�K�#p�����i}�jG��.��t�=
D�
���K���������)sF&��ϳh��^���~q�	���3����q�}�p�@[�UPPPf����\������D���o200�ʔ-3�"'�������P���p>�%M///�7TUU}��0j���e��N'|ϡ��d��¿�[�1}���@��v	����o2�=ԕ$g�ţ����gᄑ�R;���o^{�$�v%��T�DJ���6�}h8����:��7�<��؈�8�v Pꅖ�FP��钮*E>�:ύ��k��8���~��pV�Wӵ��ܱ��S�Ò��ܚ����S_�p�|[��2��/�Y����G��{���y2kx��xb����)���iӢ�������L��4�͑ۖ�7�~h�l�"�///ŝ�_d��>q�	��]����jҙ��j[Z�#X��-w�T�ۀ�&��s��"{�Do���m�Je����JU������օ|%��/r����WC^;�.�J K(��+���%����Jl��)1��������_q|zKy�Z��'nó�jl2w|w��<�,���-ǋ�b���&� �}�u��}y���c#���<��av������� �.v���ϴ�~�W~q0S>���=����k'c��߿_c�D��`Z<�Ԙ5�#q?��\snn�n`	s��n`svrx|���G�D"u��%lmm���ɳb
׃xĪ�	��u����(%��=�5�H�7U͒��˃�rv:����4Kpp(�$�����	��A�@3յ����O��@`ӕn� ��w;/�d�O�v��B�N���"�@��>~��bꍓ�#K���]K�=�w�b��}~V�ꥡ���^&4�pt�殕�nx�a��OW��:ʯ�:�$��2������i��g�d�,�>�e�b}���;���̶iY�J�^�-�
oy�!���e>�ܫ�v�9߳<��$�`k�V�?8�w��s�,���џ�'l�Q����?[���s�����{yM�	jW��d��R� �'���f�.����_��W���Z�5�\��OZ�����L�,�{�\�$y>0z��+x�ɪ���v��������`��`Y������S�5�ĚKK�(��R��{�G���3�v�:��`��7وSb��e!w�Z�V���O�{�lư[�沣���+d5��t�����/8H4v��T�E�	�+����/<rv騛D��mq����$8������ۑ􂝋�C33�11�m{��S���Z-�%j���⚛5�_�{xT���<�Y4ܫC�(P� YH6c��{�~k�.�����`#"���w�x�zw&�**�lS�o &�Iy�[�?���%{]u�r�j7j����q���-��y�񍏖�������%�&o16��Ck}@^�O;3���>��/@q�$	iA;�k����������4�ާ q��n3T¦��ۋ��$S��b�K����̪W�TGB�2�v,��oz��-�S�.=�?������H0j������O��Ĭ��s�]�㝹�o�W�n�R�؄� ǈ�zp� ���Q.����3��E����rvB��/-�����M��)©Ԇ����}r�>�'8��t%GI@�2ܒ�V��CR���ٷ��A�+�6�"�(1@|����|�����O��� q�ж���iFpI���0(�9=�?�  ���!�j�`�,R^4��``b��?Qe�^ڙ�}������]�
��(���744�y��TUW;��R%x�O������d���PܒK�^RcP?��6��h�Dk���Vdb~�q��է6��6a�h��K(dٲP�x��A?����r�OS���(]_޸8�����K��DoT����l�E*���gu>�7Rڝ!�b��X����~�䄿tO>X3=����f)��v��ɹA��˙��=�t�b�c���[�c��D��D}m��V ;�r����iX�e�g؍���##�DXn,9������D���c7ww�Ǝ��[�����C��(z����/Y{�8�=m7��f�%��wܧ�@OϚvy_,貾���릲�J�RZ�{��W�KE/�뿲����G�P<etv��$��fb�V1}(���m�R �:�L	kF9[ x5�b��psE��0��.�ʍ1�ض1Qx��!�w���܋�����q/�-1�c���9{�"��������2�&qO)f�=��S�\�<�"��m��	B�pw��XYYu�l�V���t��j$��)��cr��~Lf�s��-ҕ7����K3�Þi�!h��RE�Q��H��l7:��-���Zk
_�/�����>�Ը���A������y#���Y=�}���1��B$��鄹�L��lI �'#`�ORMԍ�
J�a�ʂ���vn��vJ�F���$��J�K��/3n��֦!��J�ɣA��$�~g��㿍@y��<��Q�7�p�5!RL��7��X�Tp�׫�|�Q�n`��ϧ�[����Ɲ��P�����v�8��W9�T(3-����m\0�OT$����r�����K.'��$?����%8�����/��Tˤ��R8�-�4�9&���o�6��A{�U�S}���T��W�0�2��N����r�O�s�_���P����^!G�?�݈�t��iQ��,�Ey�
jx0�2\i�"F!���l���/]��`��#&-��`ebaA����'��q�yW���qW,�Z�Y GFn�-��Fσ��!�`���ũ����vv|	�z55O_}n7�Y�5ITΘٹ��,�y���@�l;ۧ7�o�h��l�Ȓh9�啙k��څ�q����7�7m:#Ѻ���3��Aj�H�����uC�b!'Atx}xQ���؎�]΅��eex�MG���`�38]�iv#"u�~㾔�4_�m�X���w��[���3'V�u�O��D�3�eƿ�9$sM4kx2 4F�\�>"�pF9�x�������<j��[Y��<�Fb'��Y�4�P�#����{�cc: ��a�Y�ō@2�����w	���Qs��xx��)4��aܠP���`܍'��^-f)F�9-�YI��2 ���!�s����A��98&^�j�v�3��T,�\�vy�f�[��o@��_�y�$�(��з�]k�rB���G�g�dսl�z�an��;���x�4� Z��Ms��x*�V|�썄W�/�ˌ[�5���<�{��%j�fP�?MG�v���N�bbGǗ���^p������PiR�--�)�>LKKK��c���N����)�� j�����wB}q~I�K8\R��`���9d}=#n��ή���`hr�g;9cn`� ���pD�� ��)�J�,u������S�V�Y�VR(~gu'���W%���@K��$�y����M*�?W"�g�+�*�\"6^�Y��{.m���ʟ���fLN��b<*���o��d~M�3�p�9�����o�]��L��]p=|��K�ϴ*N�~϶�<Y���7~�$�:�~V�R?;?�j`Pbrx}!�E�&��oT��s�1���0������UT/��N�x������ַ����Xs''ʶ�6V֎�Aʐ��<EvI(555�G
4�������H���4�'aU
�RK �����ݖ���=�}�N4ų~��Na6�q#v1�v�[�zҜ�u�����S�')XR����z���r��3ukx8Ť�o(��Փ8Y#zH�ɝ��wz p.���[�1��B~+A���A�Y��3����zw㿽5H�,���������cL��fmW+�{VP�8Vvv�BQ=N5O���\��֖��߿I�ɭ��4�]]��{{�m����o��wW�_;N�7���������L��C��agg^O�<� �ITT��h[;;܏FGG�lRG�g6}e��I[t�=���S��u��|�� �A<|�4&`�nM~^>�Nà)�v�/j��04u��\:!�t����Wo�6���9����!xyZW@7���֍���b��RC�&ҹ�V4���3av�� ��s/��1~���Pwd"RT�_�u�Ay�q_���,Z�����rb�9�R����w~���n���X�	uf'��f��.��/��U�����l��{�����}a`g�g���5��͍&;;����p	?y��9a�|�㮤��p>|4!�XvNNμTMUUFv���������I�0k����W�2{Bb���5�C�w��\�C����Ip#�dP�)��������27��I���Q����i8a���%�,�Ʃ�dt���B��`|{o����ob9��>����Ǔj�I*��A�M�J��� ��Y��Z�}�j�2�_�6A�w�5/A�Z��.�`����������{��k� |��1�������T����x.�e���=3�}�n�ck������^����6�mn���S� ��/3\�q�>L[v�ل61���5��ÏO���y��B����&I4����o�����Mݐs�M�`�_�:�B��~����eT�;^�%W�}-x���0������L~�N���rCc���L���b�.Z���^��b��M?j�L}�M� }l�p����F	�c���)�|��H�Ph�8Qm���	��{��g�R���L7�O���̓;u�� ����[  �����(���v��	���\�4I����V��%t[�z�Rzy�൜��ȝp ���L}|� �V��)�231��T����K�|O��n����2X�gb�R�hV��*�1ڦЃ���TZ[k��ϖ�f���b].�Y��$���I�D���'�4%r��:OF�����GY�UR�����(7��#Z���xCf�[i2�D�^!Dhy]祊2�q�@R�0���ev��v�M��x�� "4ѧ_�wc߽�"XV��Q>�9؉Vg�Y��K�r��օȿ=�+䙠n��3���h�g z<"����-Ƈ��ڰ)�*�1b��{�6bNuk2h�ޥĜ��1�I.�.@�2[�/�17�eB���S"Ω�Z�n�;�H�آ+����W��X�U��eF����+.Z�*ff��6̍T�ۅ�$�)��cܑS{��r�i�;)��y�3�Ky����BwG�����#�i�2�Cp�i� ^�\oU�r�q(�K3E{�n�?�����"�G#s��.
�g��;�
�� S�h�mV��5�ev/v�)�eP����hR���ڃ��Q��-��gRN���G��M8��Y/qGrWGYڋ����Q���iVaֱ4����^C2ˎ��A�*��"�Ww�2��-up����,L�u0+!!x�z��B��-z�^o�*4�r�R'�9o����D�g�怯�*�}�i&��[�ۄ�\�o��������3�z	ѭ_U�M�Tl���Op��F��^Z�����LU�u�5\��_,H\,St\2�d��t8�Y!�<���3����/�������~<�?���D^�Er�d0�C�h���}��o86-_SJ(W3�0������z2�f�
�R�L��c�� KjJ�w�C�EWz^g��-K�t`k���X�N�����d G����}��"��ڦT ��?]��#�+s]��Ƥ8L��#6
��'��p{)�ݎ�j�v�]��b
3)�V�O6G���O��ud8�<���gb���fa)kM���R;�mq����-�Q8�Ӕc�>d���f��a�(�I�Zv�c�^�<`���큺�W��N�Y�2Vo#��V���뭊�3��
=	?�O����a���:ϢP��y�E�.Õ�8t�>�;��1�{�-k����-6�cAq����򞎕m�*����l��Z�Ɯf�Ŷ��!x݃G�UA(��;n�"AC�����Ût��u�"3%İ�����/�'+��j[^���&��%�]��4�����^Dl�r~Uo�r�-d��)Q�����bgI��I�1�چq�g�i/���E+nK��W_ �@ɢ�̴�z� Y�}��	��n(��=��E�%rn4L�������Փ��f�.�0�G_�8���?��O>}~1Fr9v���~��A<w#=�<�l̲�݂
�9�ŐQ�a	�tzAE�x�6G�u7L	�<��o�4N�z�9k�� �Bf+k� uիUk��z�Ս��瘸��׫eKH̦?��Y>�O��c�/BpGŠIak�w>)������8b��Χ�?��ç��� ���6	a��;4YZ���ְ�ٴ������}n��EpT��R����8(u�
���<���,��Z��`����Tʇ���9��nJ��I�C>��x.�{�*�,��8�W��X$��ίmV�#Pv��c�C��z\M�5�@f�{��\ʓdr.r?�%�U��#O�����-�6�OzRT]�&�-�i�+��O�(w���vA��z�K����[����碌��I�'�Y��Fr�-�W��[1ϳ�SM�GjȦ<��̈́s�A�"�l
4K�1���S�֒�fFj[�+l���I��R��Ty6���{e��|��3�e3��-��T%�������7<3��Ŗ&o�������>'2;���
ӱ��n#Kg*���3*�kv6��E�RyWy)G]�Rj6K�Fސxh?0���?{�JҰ%�`r|�2~�lNX��G�Z��$R�i���g��ih�0d�ȓ���IOy���0M�q�F�����eȆ\&� {ɗ�ٷ�j#��p6���0w�Mn�#�z�&!�:����,
�G�;�T��_� X��i�톇QϚ�.�@p� �8|���,�Z�v=���C�St]��. ݀]�|7F(�ܣ<�2�/ ���2���w���6�Q�܉{��Ơ��g�=ρe�<d�f�,�Na�.�\J\��4�s�|I&p2��]_EQC���1E�*�����]��EIt���I�QB���i�M�O#��eRj���}
s��>���Z;DJ���0K�(K�E�L��O���\��7�`��\��
I���8�E�=0��	G�w��|kQ����i�y���ʗ
h(��h��İ[�N�@�t	�/XH��.�����h��g�z�`��U��u�$��T�q��3BK��#g�I�`��ƩǂV�)�!q@��ئ���kN��=N�x}�sr)r��K+!���&[/�p�?��6�D�)с�,�M�f�͍U%�( �`�E���+:����`4���B���������%�zUʷW�i��in��D#)N��x�h#�uFk����x8��*ulIg���/�?���� _$�L���w�d�8����S��f&F>'�|>��ǃ;$���?��N&�
drS��~,�i�٩4j�i��o(�������	��*���/�FR����k��0��-Q\Z9+�2��q����!��3];ǵ���pD��U
�7��3�T���E�����X��|��V�W����3����{�H��-�+��tڑ�EfhB���1�D�eW�ƭ'e=gH�qI�?4���>}�}>�n�Uƛ�[�����e����]��/�M�~�����fu��׾h���Y�a���jՇ O��<f�<( X�`�zs��8N!D�,�]��>c���c�����#�b�I!�(��~�C��Q��������$<dUgV�|Wʓ�qH�%��u��GX���}�ϲP�Y�>Gꃝ8����g�4�z_L뼲H���^�x�7`V�o�*Q�!�ؘB/���8 -�nXq�Eg���c�ok/�nSu2ɸ���QC��Ee����&t�&���T%;���>8$�@gAV�=o�Gj��L��g4R*(���=���Q��k��s���u����+�<WǷ캢�袿u��:/��w�A�Ѿw&���s��nCL��޷��L�m���*��P�l�^�����(�)���%����ͬ��e9LT�4ʇpH�}x�'O�u}�e�I��S��Sy�HO��d ߬,���븡j)�}�-&�V7.(�'\�x�N�>٢{8t������k��u�>��X����La�y�RZ��TQ:�A����լ��b�l�r������Ѥҵ��I-���@���K� tAAE������'��M�@ �T��ؚt�R{�9Lk���U8�j��E6G�ף�S�Ҙsa|��C���D���P{��򩓬A�-g�-'���=u�a���}�%y�XϢC��,��s)	d&ݝ\fwYD��c�a2=��Œ#x��%�c<����g����no��ӮE����;ʻ�78���W �Y��a��}�yZ���.Y�^��7A�B�HٱST+�A�QT�1v��{��
��f_�t�Y�M�P�������.S��	yF��D�LH���޷C=��\��:��0M@�f�]ǌ�XD�p��O�@B�I7�r��<u$u��[ʾ���=�>�K���)'w<�#���6�^�cΟ��������Z��?	���F��
�&l�J�ަ��<o��i�aW�Y$�a�Iԍ�%���W[wI�;��j�D��e��V�o�o��C�7+��/��R=�~P)�����^�Za�{����KE�QY�~���l%R�P�H]X�W|�88 �4K�}{}JF�Pʭ�����p}��-6�pm�[s|�e��*j�4"��� �Ir��Ii���	9�)׈�y�M`B.��gq�z&�{����f�;uP�8�=-��"W%�}I��ӛ��s��p!�hST��5�M��Y�w�3�f9D�%�z���{<������'}Hf��|Bغ��=>��R�MN��ǡ�y2�#���+�A� k�	߄`T�)��ל�?���Gi��2\b�^��{l.�S�W{�y���ԑ�Ng��Tz+�,������ץ�Iн3/Rxޠ�q�A����=�����[֕%
|\��ꤝ&N�	7�ڦ�X2�u�o+��U�/�re5����n�i-���v=<�-��j@�Z��$�&�W�4B)�����MtȹG;�e�1���3Zyo��#��$�>�^���<v~pj�&�����_�f
�**�����6�ŭ�W��lF��^<�[z�~�xU��\�c�8=��hz������͒~�p�����&�����7�]�i��zA�l��7S�`g�U��k��,���J�Z��w�	�E[I�|M��[���S
�2WiWg�d5�Z��P���۪���[Sz*�U��l�Sޣ5�$����9P����+��,�2�}�;|���wb�AdIш��S,�m��w��N��-���\���ue<���+w�I�Q{Q�%+]W���A��Qe�w�}�@�8zv=�qjG}���w��V;j���(屖uQ)������������~�"s�ș1�6���"2�Q�{�z�$�[x�I���Gg�3�����+(�l�9i���'�s���xNɎ%�3 }��{�Ǘ�RҬ��5]W�����Yz��Ӽ�q9�=����^"JwE�-�(k�%M��#in��O��!q����q�G_��E7�CXJ��6�f��ϳ�F������vG�L�wţ��Wo�xwPՈu����G�6��p������;y�*��O׽
E!�y fl��و8cN��������N�F�����>}i�WR�JZ��@4��`��xp�C==�`u��g��E�U�Q��N�|�ƅ3ޫ�xl�+`c����x8S/�UEc��9.����� ��H�fg��L�z�!��bh.kBݡQ�/⎣{����;�L<Dm.\�X�XP�#KIZz&| ���9:c����A���&G훫�2^,+X��]f���E���ހξ�N��<Ҷ���^�
�����V_��%�<��^R� 5$�,�O&D>�m�st���Y�%�`t��W�S�P{�cC�|^�Ig���k���?8
���~z�`)���J��W��R ��^l�<����)�5c����M�;fN���/�ܧ"Dw[-�?r@/*|�It@�~G��T_��v�J�4�瞗3c|�1J4�NS�[N��W��hz���_jӱ�u?�rIe���^�6�k��o�9=��j�r�ķSK64ǉS�(P�cu�Q$Z�%ŽTmR鴢2f��K9��?�!��!A���|3Su�dō�w�7�~��oz+��~y�{H�t�<+��C�����-���q$k5�O������][ge���R�Bk|#����
�:IN�쭣��ma�{��!�~VN�Th�~%-0�ƹƴ^7/c��<o�`S+��L@��W�O�P����f1r@4jI��M��E�˸\���7F\��g�s�0%��!n�piK:!�@<�*W�:�2ڲV��Z�Dh�h�G��EhV�m险�?����%������7���CG�|
�j�A,�>���yp����S�p�����.���ڌ��Bi>��C,[����F\z�n$����
W�yD�bIhz�uӵ�ۼ��w{BA	��>׻��� s��5��c����O{��L��b�ڹ w�HRs뇹{�>��1�]'A̛��O��>��=2G]o��]naO��J�ٯ�[��&��pyd���) �.~���.����s��w�˺��e"u�7JRd���������t(;���%��zc��Vn�qd;���p}���$���#M���|)9D���|�u>ҋ���$�ն�)���<i�x�_��-/�R��Y������j�_��>�g�%�u츊a��V�uUg5�hSXDZ�"��̤�����xM@;®�d��\t=���VZ6���b��9��N��/��U/GІ���#W@~��U��z+�2Z���3c��w����`�X�@q?)Y�9%*{�hY��v��+q��>��o�3�ܢR����FW��b�!#�.���꥛�*�>G+�n�~���zf����S"�Ց��ZӛnMu�2�K{���d������0��eS�JOQ��U��e����JG�|B��d�����8�ki#�V��P��/�b�y'�HX
�vq�����������?4�W87�Aj{��'��d�w��ô�;!E'���i�)nЧ�x����m��I��%��s�NR�JV5��!�����ԙ�U3�ɹ[����[�XK��I�h}�@����%��}�6�sz�_�Lc����O;�-�(�.X;�8����9x�z9�ؚ,�2�ݿ�(��ޓ�B������4����P!oE�9�\ٰ��ii�d�������!x����Y�h5C	$b���Ч���8�&��b�p�4/�h/\҃VumNR��IU�K�\.m%�V�����1'��D��I#췜qW�ʵ�j5��/�w��'0k5��E��8zd�Oa��x� ۍg?�yI�"y�u�,���O~VV����`R�,��l��f�f�mo@���"�����l�p���_�|D�[R�4�ɨ��� |Ơ[% ��C�>GP�@=ݖ4�}�n�U_Hq���,��/�e.t�������:D�����d�$�Ąe�q�������[\����}�����k���2Jo�Df�J�ٯ���u\�=�<�����:��:n]�.88ː�8%��M�1�p��(��ϊ�Ua����=ü>����l�J4�i�7�&}�>h2}/����� ����fbd�e���ܡ��r�MHV�[>����[X'D��%��^�e���{��.U�>e��?Dy�p"�2
�B��� d�Fz,���.�TY�<ϸ;�DC���GW_J�čc�>H�Y$�$с�r
{���*P�QA�p���3���L���)����#���g�S,�y�4L�H��&7lO��HV�ũ*q����� �*&6"��$C_��R#�=nHY�}%����uB8�v� �@u������?�tB����ѺAs��f�+��^�HWj�3֏}�r�Q�E+�Dt�p8.s��q�@�c����8���x4�4qwZZ�K������)O�u~��)uL���F������� �]ze�K6���?����lw���e`�V����Њі��t�F�iq�"�_h+����:&��/��j�`ῐ����?I�P)�Պ0^�Rv�� n3X�r��o�ny�!&z��|����M�*�|��m��V�[�q#��|� 1��#���Xc���ms!��h�<>�* �:C^�)S����x7x����/t�KA!��	�(.6���i���ރF�9���ϳ�O���gL7��}�"u�'�[Ѝ�Lb�E�[�k64��?���O�j#����roX��$��o�M�㱯�w��r�H���T%p}bD�VO een������O/Y&�nr��?뎸�D��΅0�{�o�㰬_	U�Ǖ�p�ӄ�R����w�{A�ܶ��)E���jE��j�����x�ӒR�K��6��3p��*��̫�e:��\�[��3��T�bz����[�%����C|íO
�Qϐ�����b0����\2���(Y���<#>�V�8Y$��X��E����N�`�� fy�4u�x�<*��y� �!H�2�ϧ�'�W�����C�N]v)DԮg�ٙ�ѧrSN�QlfI\�"Hy�<�|��G�;����	����ra�-\�����J�S�Zw��;���-��m,xZt�`�3�ɴcJ��]��5lF=(������ʧT�R��������;�ex�
�"GO�Ai֬^�R����R���	�90�и����4���Ad#�P�Km�~ �JfXF��!)(<Uhg��P�L�ڍ�Q�kWŇ���[���N.�v3��\`.Ckn��R�������5C
>߹:0��wT����ϻ�0@�q5���~w���0O�d5��埅��ֺ%���9_���{@8g-O,1nS>sR�>��Ѕ�Ee �P���23}�:�|)��1�нO��h��Y�m}�I�l�`��
��E�Te��~�g�W����ꭣ���7P�iAT�Ni�����n$�A����CAJi�a�B������]��yך�X�����~�}�9�,_|�;vȔ]�ؽ��G�&�t�v��f�V���3^�����v,�r�xo=�-�i��һ��n?���B���B�H����@;�ү.�T�>�O��Ɇ�9�n�K�2f�$W+�*�>�	�fQ\=��R'�(�M�\I��η���v�h�<��Ag0+Zs֔hCXw�1b�?�@n�{�vv� <�y<i��ѺN�"+�!v��r�!���lk�p@��7�Q���E�k�=��ƿ��L@�H3ߌМO��FwH���^R��CN�#nn"�%wt�=����o@�-����}�k[�o5>�<���?|^^��H|��ap+�!K��2m҆�y�d�~M�Ē��+Ih�.d&��<��7���+�c�b���?G��]�
.���:��u�3�s�K3��q�dd$4]I���ϋo^=듹��}Hf�Y���?���H_ϗI"j�����`@Tc��񈅘3�M$�m�1��=���! �a@�u	f{��G�]�
R���}96���i���sQ B(���\�߈�LC��w0�7�u
 i�V��\�+�8mw:���揣�|�Ԟ��bXh!���k�=V�O�9���V��k�v�e����-�I���(Y��>6���,A���F^�����C��!���R�����'���'#�W�"+�ْ���b\�}$��d������VH���~S�b����iFş�4�h��Ӗd٣�69���.�gu��Z��D�ц��,�=�jrw��.��]cL��u4eY.�[�D4���K�+8`��wI����4ŉ�Y^�.�s���$
�K��o��}û�=?	a����50����"�
���$�!�����f��K�l�?�IВMm��F
��?���4�t��Z�-�d��.lP��{�ȖT4dg��{y�3������v�����o����R`�L&�˗R����/u$fj��-����Jɯ[�u�7�i� ����g��͡7Gh��.l��A�������߲�����Y#���S����(�����`d�-[�j�Nڑ�t'.��Vҹ������)qj�����pw1+�3���z�	΅��Byl��~���3\%qEw}��G���(���,Um-r>��BH��P&d�2����@�����8]��J����S���lw�/ڎ��H`�˳�^F���׆����������}�7j.�R�H���a����L	�vr�k��Jf��EJ�̱LŲMN�rjcz���)���. [��d���^R�K5�6ms��W�Mڴ����D��~�jmB7��(kBA��?�K`��a3�o� ��bC�L;���ܒ`�t��E����0�]D�n��}�{4� 7�#�a��ɩ%�T�!��!5�Pk�1"���)h����C�pZ^�Ʌ��p���d�OV'n��5ǋ�xOM^秵&��&���u�����X@�u�sg�>M�A`u������&�X]7�������I��r��U(�y����8-9�Qf�4<��-4�V�=��L)�%�]�xQw�H���i>�I��y�Ö%�$�W�u� ����`���
�����8y�{Q���҃U��<�̘;��sꁟG�tZѿ�����O��;6�0ި� !�;�wH�<�m4��.֬��nˣכ2~Jg`Y��@�ö
Kx���ϕ@�W:-�9U�{�1���_V�:��^КA?�j�=��$�/�1n��K��3oAZ*�QX�\�������/���J�����}��t
p*O�&�ҩ'���!0���H�ےc+8�NI�����;V�ms(F�S�r�R
h�m�zR�!H���~��ZJO���>�� �ݺ��Gǵ"��lgK�H~(������(���x�Gw��A����!�1J�sD��3j��IҬ߬�Q���U���r8O��z�^�{XR���Z���Zh��0��{�#�e����P�6o'	}�;�`/��j�yL�I	Y]�Ә�h0z�)�I�E�������x䤪�E�c�14!ݣ���n�p���(qU��9�56�t����"� A�w�������}iԢ-e�-���?2F����!^ǟ,�4U��j�l�M����^�S���V&:�V�D�����a����5H��~��v�H�LG,��>$?��,5e'�t2�N�/�m��@[����:��lk\lc�d�-��N�^����� [�<��Tv�w�g����Q��$�?�i��'J�0|����P&E������j.Y6��J�����^�J��Si�2���+� Ф�'��D|��ܹ��z���úN_ƛz���j�>A6x?��8��nxӺ���vH]� �Zv{����/�&�b���a���D-�3]#���xa��x(�3�X3`��Y����n(�$]8��;!Oֻk&G�)?yx�c=܎���?�C���wY������ag#�,��xz�M��&�QW?��%��6�J�]���w�\��(��`zu���{��y������Z�8�c����-R�Ӕ���ݔ��z����:�F�!g��!D`��&�!�(Ύ�F�#u|�; ��	�/VT	N�g��4&����Q��(ѕx�'2�3z�#ch�Q�䵼��J{
���w�mA Lg���I����J#��L�c�o���#�׾,k�Y�źq�{2�Ɂ�����z���>e��</ol�{� ��eq�t�|<��Un���T�Πz�*�ek�4��roa�mj9�\p�c]����2�W5Y�m���Dw�d���$|9g��]���/w��>�?�Ń�	]�V}�+�D���Ÿa���6���:�1Hl��'�h��@��3]c/eY�_���5��k���V$�(lA]��O/1-�����-�����b �<�����3��X5�:�:k�3ep�%5���}�ɿCn�S�;&9�ߡ��2�O��oi�6�����t����Gfp��.�[�gAa��s��������"o���_���F�<�>�gU�J�v"j����
,��d�*�R8=��k�6����g
N�^|���[�5&i�b=���z=���ƣ����X�$�	���_��Ҟ��I�~b�W�{p5�lK�ys"aruP�!?����l7&)6Ң����)"�=�7��47�~����\�����"��ގm����ZC7�ϖ�׿Nc�3�!7ߙ��e���9%U^_��ɊȄ�<ޔP�+�֟�o��S�g%I������3Z���GT(~�I}��?N�ؕ�R�?̚��栫ߨfwJ���Nt-����{�J{E1PCot&^���$��o�b1Y�n1������wx����==��X^��7O
«��9�b��6��V��}�n[z>Ps�`�Փ��l2P��J��
�J{n��@��q���ܛ�F��F�P��H���
~ .,�)�s���j1��n3�d�J1˖�*�匏m2�;b�f��V󟗺����h�������ˮ��
@�3���Y�dJ�$����t#DD��OmO�b��X�j��~�r.o#*�	giz7D\ra�������:�����������Z�F:U��ʊ���M�|�Ws���:�!w.g�Z�ۺ�
�1�)Sx���a��?h5F^ D���7�X]P��#)h������i�1^I0�$$4�dY��k�vp�>�Y�FLy��] j���W���>��=)y�q~GSL'�Gmqvt�st��"�C�����C���`	?�i6,�I��󛲪���A)C�I�>�
����eFW���i/̜=,�)�����fݬ��쾮�fP��F��b��#�^X��;=�M\������`2x�[�$���4�{#5A����������2�.I����2U=5�Ͽ����e�:� Q�ok'm=��n�_Z���pj�1 a�:U%}�Щ*�I��5�~UvD�5��|�'��G�
���OLrf���=�.����ZJP#X���b��Zyu ������{z��>	ʃ��ոG?L�G-Z�H)��i����AS�Ύ�d��C�G��dU�}�1B�|<��	N�+X#�&㉤��}K�� �\گ�_2��w��]~v��3��q��ӳ'k��yT�'[W[O�:r}7�� e�u�2y��/�.�l
@������.a}�]���Ao���n�4d�S;��*�4̝���>@pN���y`	���5r�O*����t�{y� hI��?i����$���D����n\`��=�2+��/g�^��n\aoi;~�_��Fd��^�	�G���ꄰ�p��Ə1ׁ����9r&��̺_1 Cﲢ��
&v�L(	@L.���%W�13���w>ZO���9��(DK���"7&�i@���ܿNys�fj�w ��(��g�rnd�R����8��:��������>�J ��Zh���h�Di��ӊ=T�7J�{��.�(jV�K$��!���`��������3"�.o�"~����ڤI���vlN���|�0Gz���R��:���w��00���@'�,���!g��ى�-�TI?�l�����s���O��0�:�F�����Ze���_+�q�K���WM,ڮ\�5�ׁ0:yå0���Vͳ�%��Gã��$qJ��x��]?��I� �^�_�+pt
!d�ͱH<����	�W{�3iRS�/uq���F��u���%��(SNJ
gB��-N���y+�}f}�zM�Pm�6S��n( �Ϣ���+�i*��g7�� U��d��(���/�=5� �WJ���kp5����K,I�+�׈s=?]�Ճ�z�q��qbF?���;��3)YpEk�p3B��ތMR{�:��d3�x�,?�����s�@���Z�aw�mwh=ȡ���!���V)���`Zntt-��Ώ5�fw>������o���4lm..6bBjQ��ܔa�9rt@�x�d��ۋ[wlOY3�l���5���7�
���h�Ǉ7�p�������r��?͹O]H8VO���vb����W-��L:�*�oT���0�,��W��ߘE,{5FF����<e#j���P��>�5.U-�������g����1���@�{ZMp���f\��d4٧���y>�J1/I_P�D�1z�����m�~j�H"N3�q�t>Q��ѕ��5b,Dkʄxy�ɓ���똌�#�ǡ���t��"�(�~տ:mxE�MH7��=����Qt��ѝ=͆2nD��QKɆ=�1�UKör�'��qJ���
8�Si����*t$o�s��:�~�֥N�S��4d�p�xD�A�|�}�W����W������':�E���FA	��o݅v����{~�K���z��#�(]�J��x�t��	e�P��~�B��BP��Y�9Hj7V��x6*g'���\����>�U�}��5����_���<v��סZs�ڂ�T)+L�AM�~PH��/�����u։�j��y�?��Pb�=0 �L ��G���k�������TsR�t�p��X0a'�}��4I��T�|ND<i�7��Fo��������|7�S�y��?)�$�mk��R�L��Z��)���z/S�o����8'X��G�6'�SQ2Ň�iy�ks�S��&���Ƌ�߈|�v�3��{p�x2�,Z�/s�8����b�Z�9!��\N��������:{�s���~��⹘6���2��&N�{T�Ē	��hV"�W�}���r�HV9Z�$�*��yֿ���� �Q�j��I{���z\��%H�Wx-�7�wLKV���4��8bQ�j�L�<J1rq�o��<�d�\_¥������i@�����#2���"��Jj���]a�%���ցB�Bȍ��K�E�%�/3�a��E���뎌�ж�ݻ/G�m.�yA����?� щFD%�]Z"�mda���P���"*$`<�� �;�9m|In;�1�{�5�&F�Ys�M[8��x¸���ސ�1��}z���s2ȶ)jcfQ:"�=�]~[��!��];���d������?��l��.�����*���H����a�����ݸ"����<�,��s��V�\���oO(�=¹��,)��J} q�2o�����>9�)�|BA^����cjW�xC(�æNAa_���md �_ZS�����|�j���d�|�(�=��6M��!_W�o��ۜ�a��@՞�׋�෠�bv�`�Q��_--#K���9\dt�j/U;j�Z3F���]�����o_E���A[�FQz=�&��[r.7�9�\kG
�A������:X�`��~����8�g� J qx���X�J�nb�_*0aU�m��3?_I����,s�I5ͼV�z;����^��3)�x��s�V��K� �Z��?I���.!b;���+�k�R"�w�jċ����	��I'L�)5ZT�0�F��=�Fy�����o'���������� �(SB���D�##�;T}��v~���P���̹��/�������U���&�J�^�ނ��?� �.q�Ʈ���>�)G[�ϻ����LGke���q����\�ӍSϔ#X�1�U�Xr�1�Fɱ�:`\nx_Va�b�̇��􊻲~��i�����!��(%>���o3#X��ʙ)���jז�����߄�[�wtg9U�}����.w'ؘ]����27w��(5�w�缀_7�U��O���h��a��m#���ϕ��̖qjG@��a�,����#���>���A�v�BO@L�dV�sl��º��q!��z�wI}����3l#$G,�8�{,�����o@8c3��A�?�����[�[�m�_n\�oJ�7�S�>��[�N=�!氏��iq��Z�%a�Vh�����&d�^�P�[��HF�%�f�cV��2��E�N���c��V6p/������l�a���[�/��a����������[	2�ka��k��f��;�j<s�E�}G�k�"sj�C��#��q�L7Ă���Ѱ���o��� ~QdC;L��w�f󏆍@ ���1r?r:AH�rCa�C;8�%�'�h�L�L����{*��o�@Dt�Ies���l�:�}�9�"�$h��t�NwRXZI���$�cv��ч����I�5͍��s9�B�~��m������O���I�Z&ݢ��v�U�Շm���[A	�0ha�8@���t��r�4�!6)g�L���bNyA�֝�/�s��^��ү|O�� ��L��*=�4t|��j* ���RxN*uŒ���}Q���봞*� ���v���mZ����v��ݦrM���U��f�1�����X'}��V��Eh��8Z��d��Q�Cf !���G�4��߷�`� ��R�{R=�FVv~7����|0Y��gEU���H$"ǡd�,��Cק(�74�b�듇+���>&7�IZ�MvZ��ڣ����������!�F�I'm�2Sﻡ��&�w�g�kL�I�����%X���װ �h~d�s�����H�מO�7*�a�?���YV�rw��8�����7i�s6�E �j��4���8fh)��Οz��׳s�p[����\�u�Pa;-���X	ZX�6	<�*C����H���U�	����-a+�A��H�@ta�E�n�ud ��z�=D]+�u���^<b�%��n�
\t�_ܛ�@�f����:���O�[9������-�m���su�B�TO .E:)�OIP+�G$S�����`/m-�I�r��'v͈��ڍ��� ��D]�Y�D� �Z�v��_P݀Y�cCr��g_�&�#L�8��'�>��A��oL?"gE�ť6q�N���9C����e�����ц?)���.���S�"��96f���;[vA�/�IF�����D8e-w��9���:����O~��ۋRL~g#��XO
0���i�y�RW��	�hV�ӭ
�:���{���}L����`��4�HI-ڭ�1[��օT�l�J�#�2�X�v�#��z���`B�6����D-���!Hi��ɧo�f1_r`�����U@j&M�YZ�nٳ
�'�3#
[���p��8E��bT�o��f��ƌJ����c}��O�Z�b�T��HK��E�8�N��ZA�&cu 2 ���FL6v)_GF$-�� ~D�8߿��~j���Ů>d�9����⮡8S<��3w�~=SK�	�.���Oe���X����oĽAb	H��x�J��;�N������)�ݢL��u�_d_�*x�(ĝ~�f���J�Ƚj^�N�,��Ci�o����S�#�f9UX�e<2�����`�طIe��.���x�x�<��L�iz��;�C7�g�ZN�Yo�0J�Ț�P���*Y���I�>:���ju���M����t�������|��)&�w:L1{.?����׃���J���S�_�j���il��c,�I)	��Ӝ@n'?Q�6��(�N�g��ACw�M�ly?�3wûQ�fT\�����h��T��O"y]�"��⫷�=�m�I��`�1e��m�oh�7�W��*�`���a�?��>��{Ya�6x�msSz̵V$�'�u?�;����w(�
(�hν�[s鶒D0pk>�2�j�[13�E�%1�qN�zU��Z5����U �)�Jg�K̳@�An��`�ޖ�:p~eX_Y�Q5��_�y���>kEn���&n!\�]��l���G�xU$��3*	����5��!��~U����q],B��n�釘�4�n����Jy�ދ�W��i�i�{%���J�[�,)0���Vꨇ��8�bi��8�JZj�O��&:��z��;��Y�)=΢�z8�\��f7��������\���'��I}�'�Ļ1����P`�7QL%v_�@{��{� -`N�G�0���}rϽ^4���q^9%M��]�q��ܓ�XHmPI����[�(�[�L�<���^�䮊ܓK�)�<�]-K]�߻Or%D1�')����:����;\�4���eS����`f/Zvx�B��N�����1!��B�5>���_�y��o~�\����^�.�SQ�JFT�M�#Cd�6����I�T���%N{S�A�4��C��rX+"@M���q�{'s�Dw_,n*`�?��-X���8�ͻ0�e��ۈ�ܖŉS��Kqq�8�j��l���
�à<�F�ԙ���pE�NP��I\�Waקt]��4��+��R��I4�勆.�����hN�8�~����Ĺ��I�4l���x���Z|��/��@#�W�q+�&U+t\�Y���� n�K5��jՐ�6gS��0�N�]"Џ�hգ��!vU;����i�*�0�9�c-�	��\�S�W��%�p�?�z,�8��Ҭ����W+���P<I��ȕ 4�,d�_�5 k��-Ε�i�@0��	"�OT�*[Si䜁G���j�	���%�AE-��Em���E��"O?hB��Q�.�虜v�` h�)~�ôፂ+�#
T�h�`eڭ��CV�h��C��,��,�����׬R���7d��%��?��q-�>�u����$��<)��G�;�8���H:�c/>,�+�減F�KUf�D�3�\q�_5�p,��/̕KL��zQ":�$�9�
ޖ��v��� ��tP��Pc���6	 ��>�k��C��2nj���N��T���B�=R,ع��r�*mRyk���q������¡�~�D�pt������c��f�k�Ϙr�/f�ݼ1qiH���6Y�sR��p�Y��R��i�k�[�֦��x)jS���"��A��DD�*�F(&ob\mW��ơ��e�3��"GkM�m�ŸMc���ڎA�Xn�˜�b�T����I��CF$$��9�q=O;�ݘ�I�4q�\����*�7v�Lb����)�N㵅$o ����� �NU�'��D���3Ȇf%
��Z4<��FȣL�n�R�J�mG��O�:��h]�5�y����ۦ�Ӡ�����^j?R9��ۍ@Gɦ�U[N@��Z��W��P\qY����O)~�FnJS��R��P��^�LƄBC�l��GSN��9b�(��=t��DJ$\7ǥ��y�����7���Uva0�vc��Ѻ�W�ō|���@2���Xe�h2�:ǄBbd��%ic�tZWZ��J
���ƛ�~mM)K^<��_N�jζ�_gn?y�,�$�.��dW/^�1�݉ީB��l�;���k�`٪
+���>9����O"�G�0&�5I���Gm�t4���l��"��v4��_����'T8���":�v�C��O�B�R���L6o�c��r�z�ދ��S,��'�}Wҏ'��Q�g��{I���b��t �k|�u�AS��|�_݆��_��6x�g���$����[_�kG[���i��Gw�1��\��J��K�<��*�S������R�N����z�Q��)LE���(T��~�$����G�
K�lN8����=_���|�"���ϬW���9E���2���|4Ԭ�9��ؙ~�OK�*K��F�B�D�("���T�iI#��?U�	�ԛ��w���̽]_��t`�x��^c`I�g��IK)E�L���
qA�)���]��\-�ϕ��g�Z։�\r�PM��Y7�Y�C,B���� 9	:�dϦ����9b��z��D��B2�_ўK�ܥ���D��	9�]��|h`/�}�{����T�={�9-<���%����X̽��1����|�ʅ���y޽ir�.� �цh�=�+�ɲ��^%@E���r���a�zs�wT�����͖f�;����}��c���XFt(F;p�$'`������Q���Nbt��#���Z��ױ�􎀝�\��Tk���}��'U�c	:G0W1��Z��W_ �QCU���S��E��o�#*Tæ��9�ϫv���R�ߛ�?�.����
Xǒ����-N�Q����P����\�	�r�`H�:T�v��R��'%F�iX��⽿����0}�ӗkH�#�$����4��?����͉�CF��;F];�~'��_�Zo)NG��i4]��]�ݿK��T����c� )E@��Dc�o��-�,ؕOIH" �~�;���� �7��v����h�{H?|�������6	�6�6cR$���*6D­H�ѐnŒnoBf+�2���'�&�s:Უ�%/v�}k��?�d�n�AD�O�n��̻	W:,���kY�>��k��Щʕ"�Nt�Mf���t�,�B�����0�_��k����%Xw=�o
��ί�:F�iHhTjIY�j�P�V��D�7�����}��i7��$	��A����Q}:�ɘ�Ǆ~)��dDkv�0a�?VĨ��"c
�;Q����֍��hːq��"q�:�f������m�]��(�븤�F���u��e|zx����Ӑ��;8��7�i~#Ɇ`��A��E���*Ro"���2]l�6�u��q��L�_`Σ��>��*n/,}���(Esp���w篾Ҧ�������)08�ײ������[o�b8�4^Z,�a��lP��	 ��\"�×�ĥM�hZm����,A۰mT�����4�`���E)�q�!Nr��F��0;�ٿ~}0p�8��?M�\\��X�DW��>����W�JN��*CQ��w���&k��u�`�B�L�{�����Z5���k��R��%�ũka�(�@p��A8^�%f���B�G�Q�����9��-i������>!7%j{AG�S1B�b���&��� ���|�<�]&+�7����}EF��GI�G�z�M�����V'dj�Xi�,�C�޵�˿��ތ�;߻��z	B9d:�Z!G�/��]-�\��&�xZ��F�a�H�_m2'81x��
���V�חJmp��5lI��T��\>�R}��9�c���YF���K%o��}��f)sR�u,ϒ�I9��O������ �2�8w�ܺ���~�v�`N�x�̩��^��Ǜ��|��7U��c{���O��4(-M����t����!�Q��,ȓlɞ6��qTe2Sbo65d��xC��Z�˱]K�+x��P�m�"�zF�����B+��[��k��
W�SBc��*�"�9M(M��X,#F�n *%5J� �Z :�}��7���B�UȲ�*X2%β]��b�� h���<����]3�@{˦��G��<U�&�h���p
�9c�{ڔ_����2�l6�%\EQ��3�D�J��G!����S��b��D�/ �7��3~���o��ܒ~��Ö�W�f���Ty�1� �0��B�9��R�ϔn� �sY�r�mB����gՐ ;�㍖�ΎJ����Ű���p��3��oķ��l��שk�m�J����Gof��y�l�a��מ��톖 Ŀ������g����ҷQ��&�����-�귋��+Q�gD@j`������M��<U���S+������Fj[{���G�5�o�%��ۿK�*C�$�)�Y��#V'F��A�Y ���F�%|����47)rq����j�E�\<�@V����Uh�ށ��V��Q��O��V�]��ɵ~��ܤ��3"t	��٠>׹.�qJL������|�}-����a^5��M꡵�����Ӣ��u���� /�t��'߆���Vd�zX�Aa���B����(v��=�tkuق���?�p�;���imWN�y�4(,\j�'���f�f����c�L�ɂ7�
^X�^�4�`�Avp��DF����헁���7�� ���1�>(\�ݹa�r=q���v ~3��w�&��R?K��8m\���V~c���z?��s��='
��M�_�6�;��R=��l���Oq�;�eͿߕҠ��	08��q	aR2��e�f���G�"Z�ӂ=���yfO�����%��)Ac������ʮ�������, ��9�r��I %ՠ&�O�3���Ј��'"�hco��i\�4��G�z�ZN�ݯ'(���;^�1|+�`���%����b!��Fj�SL�;���*����	�����7SNI�G�]�����bLm�IԖ<��S�S��J�ޑ����ם���mf�2�eCGA5}����g�Tk��ױ���ۻL(��*����[t[-좬�R3�:HCE8�[k��"T��2r��u{��ć��)��q�3���B]�s[����x��-���M�o�p�HH�n�o�s��ki]���՝:�x����U�谥z���%�K1o|�u}@��t��/��-�,5�A�Gѧۖ4�C����
tW�N��9�јA fo��C����:rqkNe�g���o^(1���D�cˤ�W�;�.gJ�"c�q�G�h(\n�B�Vo�.Jپ��G�]kCv�B�Ă�H�'!pGJ��d�����z\�QpK��JНᤙ��Jug�:������c�XI�UӰ	�[���e,0��!<45 �Nq���1����,����6� �"�J��V�IX��Q���)�G�ֶzz|��*:�� �aɀ�:���p/�'�I��j�$���t6U"����p"�G=cl3��܏�>\�!�n��w�o&=#ylG�n���Xw�%@(�PX�K�d_S��7ίv2ʿ���%�Hq� ���s�zɿ���9o��_�#%z\%I>W��ZF(����j�=m�K9+bM�F���,�}WhƎ(W��% x�Y��0�)���$�z����_�-��_������c�w��l-�Id���zp�n�'��k `��x�@�ߘ0��(B~i��(�j��WȔkN�4��"`ɢ!B� $i��Ì;@�����!\�|g���b��U��.O��u��+���N�Ԡ���|�u
�y���M4>M�ʆ�d�v�~�G���`h��H��p<�t?�	J�N,Bz=6��W��TqH�`~|��@�FWa�w�OS�D�	��4�4f0i�-+�f�\���RӲ])Q+�k�`�+	��>7��Z��X}�i1���˧�DbS�ʛ���_��W�(N�S�߱���%-�Q�d�ŪW�:�Zhg	������7֟��@�
�Yp~�DЕjP�׬XZ��>�z�f�zW��E`��Ί���y�����::t���p0Ư=DpH���%:��}�s���9Avh���L�a+��ٮ6n7WC� 3%��~E.�t2��\��2�� ׺G�ّA��4�����.�c�g������n!���]3N-�<W�~~&(����p��2(�0�գ~;خ5Y*�j7�ok0�6�����$�XJ� 2�y�Ibj�n�H�r�N	aO!���QV���=�Hr�t^�Qu�:�M���ӧ$�HZ��{N�]n�x	��"^xC�|��+��O�z]\}�	����?��OS`d�x:?�����d7Ͳ�,��]97E��n���C��C��:wcF9�u�hi��z؋*YK:hi1f%��ز�-��R��h*{iW"A{n��豚����xo���sRSק���5���rI��H�
�ƕ�[�zu]�W�c�\�J�/B��%�q��[�B�̗��z�X,,͛�*����ii�8����Ģ^��j�q��B.�`�1��!�۴%RT��Ê��2 ��~��KC�#��\��I<����Y���E?y��[	uX�T�.�?�3�Q����Ǆ����q9I%��5�f^�όS���M��DQ�]_T�iS��P�̷��j���WsM�5
��4�u��8󇘽�]����*iC�.��=��k.ب���Iy���:�ߠ��ݡQ�y���c���%
O5b�\�׀��/�jۍ�%�y�ߩ�a��i���S�]���Q�<@b�LC���x��I9��|�:�a~ʰ��;u�s����R`]^���PSJ�x@�������m��s�O$
+8��A��4�`��@���ʙ��ظK�s�5�Rn$�n����h~�kdУ����{��~�!3%�2!�o&��FV_ns Z������!���c����'M���� �Oh�~n,�a;_g�Z��r��Gp��oA��%#��� �~��Z����&K�;��֮쵑 S��]�y�uc��i�ӈ|�;m����j*T�z�U�2���<-H����im	1�:�g�"1Yr)Ӏ��1�-2�_)� �-E�U!O7zY.^w�/)K<����Y�]ٌ.M�F.� v��u�ѓ�[7�]�3��kɓ��u�+
c���/kq6��
����Z��;-%@�.��	Q�ֹ۠W_�!Zd�l?F;i�ƹy�U���Nb���2�_+7��}g�fp�����+p���){�f��:�Z���eX�]��|!7�(�����+�+lC�&5�y�Y0|G�X)v���v �]N��៱�(����~ƃ�Qf�A���2��)A��,��Ja��^��7i��	�)-�?9`v��'�7띾���RŊ���c�����Ԑ��}@������pj�����{x1�Y0�D1�y��):ç��d��q_Dfh�d+�^Yh�/g��A�u!2�r�M��y�V#���>�0��m����ѽ����-&�u���*��x��I�jB(Xܚ����n;dQp��sH�&����#(U��v\�4	���m���1~0��v��hw��XhN��ş��"/�_r��u/�Ē�3��b��EgM�a��dM�2,���i��X�G^B���ޝ0!Ԏ�Gz~�z�'�M�Q�D�}2�J�#FUf�80��?�xa$�~�~V).@ ��dJ����<ٶ�L�������h�{]������s��R7��쭃��pU>�ĭ�>b��1pT#^Z�EYZ9�O��y��>�{r��<s)A�q�%/M�X?B��!��3>�&�Ls���h�?�H�Cؽ���%��e_��-��!����A�7� 3�-�]Hoo���BkQ�1���S_=�(�5���g��K�2�K��ՂQ�x\��.f>��+m����wG,�/���Ŕ7_V��31�3�Ũ�*��W�5l�{�N����b����i���H%���j�e%>zز+|�f"��w��r)T��p��'2%h�74(f�_��n����J�ѕٞ<{��"��I�f���E.��fp���g������t�^J����6�a+{t|�8h_[��S.}�����7EKV�p��絯N!,Ӻ�wñ�ݕ�U�˪��3�����}��O�^��@�*L?�~�j7�����(�:���%�Y�L|vf�F.����Q�eƪ?�=+����TP�`S�\=�P���J|'��mN� ��[A.A�X�(����;��[<X������x�\���*Au��"� 4�~�16	yE�#'��:�7#�O�C��W?x����<+��f;�����S�jif�/�
��S�z	׸8ÿ�֏d�c"hɞ�ڢ��+
.��.~��NR7�z���Z�}8%bɸ����u�s��(��Ά����ej��t��/ ��ҫ��2^�(�b��^�q-�tc�P�!:O��r�@�zG��ؙ��3�~䃒zp��:&)@�[��:�LS����{����TȇEe,�Ą�w��)}������/��͟~���������}�:S��J}���$*��F�J��?d�T�]�-LKq���S�]
�P�ݡ8���-�Z�]����Z܃��~���ެ�E��9{�����<	���`� u]v5Jh���m���"Y�Y�ra��(:��d�$Ƚ	�5�7�D��M/6�x���2@���zcj���K����G)�/Ǎ�*y��#.rȲ~��S�;ώ�9��ʼ���K��@1.sD���3-(��o��`c�DА{�?d��ۯ��	"��6��-�"
;8��=Q}�^'$&�HV)���eF]d�>��������Zm�*��B��~��F�Y�9a{~��Z�������P y��8���(��MPg�D�NC>j�80�.�@cQ�^���'����4�Z,�
*�kѥ�օ���9>_�\������m*����j ��m�c��#Ǐ4w��?����N˴4q��o�\�E�Wll�jG?	7�w�"Y�w��Qَ�I�[�f\f�Ϟi�=��g�u㐈���{���f65�~�	;<�V���w��������d[&Z�ߐƔQU��4#�(-��C���4�$��j��B�Y�8���4�� s�����+o��~��W:?t�������i>�&�c�/����e?Wϴ��~=�ǝ��NbS�G����g,�~1�v���H�ڡ� �vMG`�[)����q�+��7�����Nk:��j0�5����e�G\��Z�h,ߒt��]�(F��"�y��q��V��L' �!��d�.�����3K��� 3� k�%ȣ����ꉛ<��Ȓ�⊝��>�IRO�r�<g#c�-?��P4���Y���M�9������]��l\�Ÿ,��V�x�zHL�E^�~+����B,b#䌃&�1��Y�b�E�w��y������rLxU�%k�O��*�뒄�'�MfJ��h��Or|����Y��m	^��Y����Lu8��)q3}\ߦ[V���Þ�<����a�W�5�f�sVZ�$��ݹ�CZ��w(���W1������x� ��7AT�rlT����0�q��D�P"|u�~
P�ʻ@�6�q��o��J�H��p���k�C�v���5 ���s⢤@��)\��u-���O��H�[��SϠ�Zr�!u���xH��AV	^G����!j�ԃ(!C��l����w���:��o�y s�u}���\Hһ� Qi����sѵ��y�3���)^�g�o�/�B��4�W]�����$@N[�DsW�"�
CZ��r� $)��L�<R܊���~fƴ��AK��������:��[�}��`~�4����/s��-�����40y���W������2|���Uꬌ�G�:H]$G9�Y	���W(6����59�������G����j r��a�9&�_��W�-p���-	 ���X��[����7�/QZ�����%}F�����UW���Ţ�@uڤ��v�I�^q����V-�Br����F^`l8?����(e^4��d꙼���[�h�ɡ\�����y��]"|W+����c]�8�O[J��K_�梿��߬�?�BS����mty�AR���!�d���p*���0��-I�o��uJ!�0g��n�?-
Oz 9V}zy�CD`'��ܹ�@D/�����&�u������Q�]
Z�8��#%���ܬC�VI
$n�`U�X6�M���Qx��R�ʗL�d�̻��+=�񰳤?5��K=%����IR�Q
� *W�U�>%Ѣ!��%w�)�-З2O����]00ϕ�����P8��F?�EDEX��\�>S�+���wq�^���{�pё���٠��'�S���IĞJ��ZȜ_ix������b`���Jv>:R����P�axUJ��Gc��H�4�hiE/W�������C�[�25=A9G�^BF��/~GC���c��l[����r�|`H|y�c��h���T�ʹK�:8cM�;���5)��q%�9���3b��y��y����O�2�<�6�������=�{i���f�Thm!�9ou#�Kv�E;XQ�K�aEw�nS�K��Bv7��[��6o��.{	]L���<�|Ѳ�[��)D����뷣�	��Mn���n%���*���~%gQ��},'rƶ4S.���Y�͞�[񳙗hHV+Dh�ЫΡ���x'��(��.�'��Or��a@�[�NRiI�aJ��tȂʓ����;A�<��^+�1��A�[� ���H��#D�|��%�/Cl���.�� 
�n�5���{+!�����&mA�~����
��M���a��A�o-<۹J-�
�YҖ�� ��zg%�TAp�����s'x�R<h�5l��N�3H�L���Td�R�4���˛�J��o���`��V�;E�;^�b�������ؑ���-�/"�ɱ<[��v����I�8� 1�[�&a���xS���M�ŉ��OG��TiE?!1���x���0���E�j���nR�RC35J��� �Ț�-d��;�>z���~S��c�}r�iu>a?����vo�&j��~��AÖ<W��s�_4�S��6�q���n�L��H�^V�jq�#?ycW���MƵ6T"�:,N<�^~]�e���z�J�����A[ ��لqozt�W{�_@\ ��i�^Юn��N���dwoA�����8K����&d5�Jz�oLk��F�HS�zr4����4�m��4)��Z�}r��'ѱ����_'T�^�YO�ep6��r��{��Q����|�H�NE�P��q,5]|�娂��I��8<��x�X��Q�%c=���� ���h�le=�n�S���iEp�y��p�?G�yZ���[63�vy��M;�`�z��V�d�S$Ym^�W�.����AZb�;�h�k��Ԡ��M��O���L�n	��#\ӭg�t��$�����97��Pxę"�o��v�+?� Ь*1���tYZ^���
�]�����;u�Ǯ��`aAЇ��kz��.�+2���ӄ��޻
�G�9͠��8���7��|�F���QO�0�t=��ס4��.���x����]W
�%1<��F���=��ϋ�y���5�7������+ZS=���h�X�F�<<�%��f���[w-������K�Q(���e�NK���h�u�O��G�Ztg�-R�,R�Ń���ɴ�ʜ��Jw���bsީ*цN0��/K�kN}�
��l>�Sgm�т.u�`��5�W�BM7���Փ�|n�,YZ�&��8:r�qpbIX��V��F���6��O�z;+}"��ž���	ͅ���LћV��@wu:�$�4���[��}�f�D�w��ꆖ���zF'v=7� ��e^��)A�uX�v]��Y9�ڼ�� -�t������sK竬m�aq5놪V� 6� �2b��RaI:��_o_�jW.��1�A���U�Q8�*�P��Gw���[�����w��<����)ƉWJ0k�ׯ���{IB�g� ��hgQDY�13�A����uʛ�X�e�O���W�����8�F��c(���h/g5��e����3e�H@�Tcҧ���ע�����`�JV"V��E���9���>X�Y�4S}�A�0�_h���1�)��t�[:�o�K�)�bp��&2�g|n\�VW��b���B'�KX[{�Y?t��`��zǵm���|<��Ӓ5�r/#��6Я�e�!xÕ���x�	cFef�?_�y�u��?��O�l�#�-e��� s�Џ�v��=ז�Q����T���]���H]�,�Ǯ~?���>d��
J��\�o~��hp'L
W�
��[ ��v�ť�"S��\ -�9��� �N�^ςRn��3Y��`�02�`ba���,�1��V�����к�7m%ɹ�Ի�w߱��xH�����S����"_!�)�z%�5�#���Y��l�=�3�nz�jL� D�}\X�ˌ{Y�D�+����h��8Fy��������'��լ�g4Xs�������c2�����b����z�V��@�T�?�LW�´���v/y<���G�y�=\����\�,VC���J*\���[r碫�O��"���^B��t��D"��9Ok���ɟ%V�{�*?|}�P��;���;v'���
��T��_p0GvI�z�8N]d4����뎶�J=��66j<���:.�]�]�5�8#F"M.>� *�,L�7�;FԸ��=�&$���&a�9:�;��h&��%]��B����$$����jv\��F�J'��"Ύ�����%��k�uo�)���c�g9��p׀�S�z8e�Q4l�z��>�|���pl���B�� g��i�K�Z�%�у���y�zj0����;��͇�F��u|� -�΢m�c�ݬc�Aү��5-!������Y��lӚ}��{�aE�BC��ۯ�`Z�g�ou�+�=g9v��<V�l�Eg\�ܟ������g�q��X%=P.���_����o�`�+��Ɩ�%�ሥ��F6������V[��l��nI.T��2R��U�^�eObZ���N�|�5��e���i�m��W�g�W0�*�¥x���֎o�����NY���ك/�`@>c�uc��-x|Z�F{TX��VeS�.p.���R��}0��H�L�	���n ǌ�x`�ap����%�=x]�ٕ L�x:}�+a��4m5ˢ�ÓV�=��P���
�bS�]
X�DnU�0���9�r�L����Fol<�d�[<J!��}�I��0�����g��i�{}����ϵ� �4s ��~#x�|B��v�}�����8��#�k��	�%�Fy�j�-R��T��&�KZ�t��0�����P"��kTi0ź�Ǉ8��R1�� @$�[�n8����_�C��A5g��9d�X�z�E�P�!!�{3&&p;G���.q��̑��,��q���r��R�8{b��!DȍH�i���n���#�D��L#������k)�ȵ�����#Yt�6߈�<tH4�K�ƥY��cv����vy27���\�B�&G�N$���i�/-���u��{��U�~]���U�YYl[�t��Z��|n��2u��n.�p=�6u�tR��b�ݐ��~9���B�XB���l˕
��c�4�8~;gT�S�ծ��V﷐����7�녵��F?�Bc�2=N�s��&kv6(�Nɴ���>q}����Jf�:~R�D��IX*�����/��j������f"�J8p2�\q�l��)��D��;HÌ��@��9�f�0�;`֨��o�ʁ�~"c]|��\[9��U�B��v�GǪw��?
���3�or�!L}��X"᷺�
��ȑ�ᑽ�x\��N.����fU�(;�u�M�5��ɱ"O� ��� �nHW�5d		�M�)ROC��H�k=�N]l� *���!�f�+��P>Z����RyGj۳ż��GL)'���=�{т?�ڜf�{霛y#۟�Ei�m�Y��-x���	��K���l���I;���F�;6�����������Sw[���E�X+��I_�{
״����e�:
_gAa�ʴ����^�ŅC
��;�7������� �?@�r!�]?}Ü���Z��{�sӖYJ$����R����l%���6�T�o��������#��n2���C��X�U���w�A�@�k`ےі�3�����8�:[�~��5#���j1�@�y2����f��<:���:!���K��=�L��t�$��_�;���S��\�w
��mh�h'���k@K�
y猲k{��-R�0�L#���
�RT��إ����Zx1���W���0�s��{��`h��G�V���� �����K#F����}�d"���Ƿ��+�#5�jp�FO��ij�D?#�I�TZjDmӏ雛љ7.OsR�2��36ZN;���������4|���Ѓ�T	e��`a�OX%�%{!��H���ݘ�VP 4�C4*b
pvv��!�6��HJ�k�ކ۷�a������.n��<�LMp b"���xI�4jn5|	g�)����W;û�� ��nf���Z�JZ=��� ��Ot��C	#�Y +� ˨:WA�\ �)1��ZЊL�;�[P��/"���,ū묽��Yo�F2�?��6���ـlސ��t��M�:�'���y�'Q����z�X�]׶���� ��*�����S�KN� 7�'u�{H�֪<��*sXf!mw�M��{�������[]o���ĩ�d�5o#�!��4W7,�s=~c����a��$�2[�]�~�Gn$Y�wi[o��T<�ʵ2'��h��ZW����\���.�XW��+RG�Sʾj��Y��'`����e
MS	���Q�'�i��S�Ê�X�L#�yg��(n,O�V��(X�X��F�M����JRd[�E�i�V�i<�>�8�Cz^g���ml��ث�jm�Omtp���
=�=��h��C�m�鐔�C?�]`�> $e� ��*��x��Ar�W�j*�."=�k��Gg�#U��
a��Rn������YH��M��2�m�|����E�Ғ�7�V�ңL�@�}���O� ��q+�ΣUݯ�L¦��{[�}��U�n���}�Z�s�l�t�x�yb"{.쬵�Sʋ�]��I���0
��#�����̡�q�<!F5��8����AH�֞�ۤ,ިiX��Qy�v�m6��̀:#�l��L����$��q�9��
�ء��EZQx�<c�L�g��=D����|�l�3�R��H&,�vP��U�#ױxU��݅�9�%� �f5P��p�B�\b�>�@�cɩ�X;<��w*b�����,��P�_�D�hU^4�I�y��F۱ǣ�='�%��Z�m��K������ÝЊ�C�ԟK�Y�<����艴 ��Ⱦs��D�W�d	�#����Ǿ
ܫ)Xs=�8����J��9*8��M�D��DB�*Q��f���?�˜A�eg~�4~�Rӯ� ��b��������]����o�g ���P����L�kX)�Bs��ҖM�@�o�=�h*�x��Bce�ύ�j�-ݿ���e��LU���ڢ;��������v@�cLܜ��v�S=�������f3����:m�{ߨ^ƣ�0\3�dZ��<\t�v���p/�"��P&ɘHH�s$Ij��5��9Ue(C��kM ��paVA�g�)�����w�و�+R>Mfl���NHO����v	I�n�J���+z9������~�����3�%��,�O֚��ñ���g��L�>��]5;�`җoJ����h��ҩ�Vk��D�L�P7�{ϋ�i�n���t�P��ί��?�+�������h߳'G�V)}���?���'-JW���yDR�7�ɦU��˰dbd�����#�8?�-�}.3�y3�m��d�s!�~�6!�{ϼ<*���H�r폆{���P�~��3����"����H��yՎ=}Լ� O���YB�����ϸ�&�g�(\�����6?O&�apMM�*|�1_.>(h4~��0@2r��l��h� ���ǹ��^M��`�a�ڜUv����{]H��(ה"�:w̲b��~�уmD��&�]�/���_�c��{?����:p�嫻`��~�t��SCv�"Ay��n�CA�q	c��K�ʍ�w�������B-�sI�qij��!�AZY��ݼj��܍<���XL�}4�i��G�\�F*ٚ�r��)�Еv�HW��t�(Yiw7�]����V�l^ʼ�kh����sN.
��d�u;��:����a�_M��mH���w��I)�����Yx�#��!��x!��������Oc֣{���E<��F/��^f��т��nU<iKyZF�w,�.ey_D��<�<u�0��o���b���s��Q�;���j^D�v��/�78)`�� ��h�ŏ�܍5��}4mq�TFg����1lfI52��]���J<�]O�h�X�B=�5ʪEx���<c��Y��;�6O&<����-��d��P���[c��:Yͽ�b$�z ��'�&��z�
q�����֭/	�78x�p��5*H8;4yX!���H�|X�}�cg��&g=
T7�1;�)>ݰT�\�I1��hZ Hh:ހ��a�m�l�8K#�p�x��:���C�Uy�J�� ��`���O�ΣfF�E7��NᛦW�
�~v7Q��G�LM��B��}{���U���2z�u� ?`��Og���gp��M��ώ��Eg*u0����a��(���\�u�	���	x#v�;g.:&�����a�03"���BX�����S$�F��k������-�cF�N�C��5Doy=?}������RRi��Y�Z�u� 	B��� םa@�Ml�n�LxJ�1m9�^TQp<ޢ+��jcm���`1A=��?�y�VQ��|�3��|^`��}�Td���:]&0���W�
�h C��ib�9F��X�7�¿�_(�F�=۰�[R��L;�ڼ�nC�wo�#��#��ݴ6��f���QN��M��zr��V�:��)��!�ÍD-������$�6�/�$�K<�l���:��[,���nz�~��i��Er�R�b�z��I�sFٮ�54��2���8�#�[��K	��M��%��=�b|�z�-�J�1Q��F��=U[v�8��9�zY�����t��V`/�^�W��7��ӏ&����k7i��>�T�?�I3k�^�p*���+(�$=g��9Y���c=��~�[z�U��x�d�I2��B�~��y��匓M�GFA`d.��t��:�
�s��k���v��gA�Iw��M����z��w�ܴ������'>W���5�kA�NĲ�{؈�v��c����]Gm�BE���.	�B��,Q}��ܽT>*r�BǨ!��7��u��{���'s�A<Gn�״�R��D���_L�G��y�;	eD��)��uB+1
����CcR����O�PK�7L�k��Db��� ���  H �	��ms�i+B�Sܺ�G4�Z��^Kh��D{����G�Ʋ�ݙ�ŭ3:���Y�'��Ì�`zA �>rsR,�[��������U�C�͡��i���M⟓�Ք4��X�f┻��?l�R`4�C�l12��"4�g�� �H�Yz|��k��zۮV���U�B�/�-��jPa�Ң��:�4�@��?�3C1�}�ԛlnT�L���$�|�c�ѱ��Ħ��(��
ۭVa�ed>K�O�}|���]N.n�π���^�u��m'_�@æv$�~6K�W�|؄�k���=zm�0��e�5�I)z��>]�B<u�5>g%��k.O׫��<��h\�Vn[$�\��ӣ3zO��O9�\H^n<0�����
Z�	Z�d�����o��-�py���7'q����'�O$K�RS�對�Z�0zP����Ąx͗�����5v����t���f}9F��p�t�
�)d�s���t��tqW:�g��pl����B����e|LMH��N9�1���Xd�B�l���x�Y��1G\�� �꿚��R��&���G\~}���P�\�3�@%���l�����p0�t���hZǗ�����G8b��C<�0>0�'�k��Y��'�CU�Qa��O>��|����o���M=l:^���g|M�!*��6�9��OI�%������
�?cqȐ(������o���d]o<�h��V���6=�X�1�>6^��&�{������i�*	��T�`]������������}̞���eR-�@�Y&C�{v�+�_�\#��P�Xji��m��W�V+s�6r^sW.:�kN�<��z6h�o��D�}�X�W�,�ƥfz�]�;�t)��rI�!��DI�}y�m���H(�W�{85���M�kw����=[�������w�t�dI�517��*T�!��&E��O
�Oi�d�d��������D1_ƙ���w�~"�@�y<_�w�	lw��C�yko��ޑ����o3��>��G�G=�Q�q������i�V-|�Y��Y�(ՠ�QE�8�L��f��j��zy�5������'|�)����Mv�~�C�x˒#6Z���A(�ۿ���nYs:Ʒ?�<��=�������?�::�@��Q����D�r(ֆ3b	�H�m����-i��yտ��z��ҳ�[C�f˚�3h�I� ���)��@b\P�1&�$�V��{�v���S��g/·���'��@�C/����������n&�Z�Ów.=��>g��@�R��E]��n�(#N�=' �𦇪-�3�U���ߗ��E��@w|���2���y
��|�qwF�hݨN�����OR۹L��o?J3�h���r����}�j�z��QW�}bF20������/��jI}m;�s ���z��8�����񷕞r�|�#3�0�X���@A��`I�kQL�-�����q��FPqZ~"JUGm��R���x��G��������T�=U��o�E�~�]{%�c0�C2K�7�C��=���;r����[��p��_Р�F�ƒ�o���6�-�N߼������N	�%����5���bBˤ-��.�m��_�RM��1����r[ۆ-���RJ�U�*f;�_,��7ͼr��� �i�nON��t;�Ϙ��f+��3���|�_�2����D��D��
K�� Ōg�Mѩ/�ZOs��|+����cy[H��|�����'+g�:{��!�{���w��̧�O�ZV�8%o�q�B8� �D?����l�(�K"œ���(d� �s��4zT��v�b��CPm��9.�:��ox0��u�F�+��/��׺�<�e��g�'��7�OE�	�u�>�.��\Ԝ�<[�c�ƺ�P���0N����7�2�e6{�m�����@�� ���2��t�+�\S6���E�����g�C�9�\���!ӭ��.R�Q�Ё�{�\��C���$��y��b$���>�y
C% �̩��8�g/{��+޽��m�a¯j��{�O����2D�21�p��|R�j�C������V�\
�ot�98��e �]�puC��#s�`���
*�l����r>D��͆ �f��P�\��&�k��&��]zb(�wzXp����Aْ�,���$#�*Z��B����7]t�Ǹj>Z��[�sJa���-��9Gp���uWC9�+��R¯^
5NJ@��7o�A	�n`�e����֣y�N�<��=�����菓�8#GB;��]k��G��̟�9���87R����'��Cn�����Yʀ@�X~.b����q_�}Jk���QKs!gG���2�b���D�����	���.�h�xo��s���]�u�@k�h��t�B��ѩP���WX;Q��Ȓ)I���9#yɴ�mka�us�d�ϧ���`�2-�K�'��N����T<ש����H��M�:�?&�z��|��ם�4�S��d~���d��L�I�]���V�U�9?�Cuk�Qk���b�c�%��o6W�J�o�3yC�^��Wn��^�̘�Cfq����5�}&ts�S�}��Q��9~�|��Єt�@G�ĥ��5O���,~	CUs1[9�������C�/��?���GݍV�������GK*`5]�#=_˺M���kY�\����tN���	�m
�\�x,V(����~�}#j�t�q�@C[nM"NoG���֔&q(�q�ܹ
����"�_����۸%��wfvT�[���űl�/.>���Y �u�m�����뇃�G���p7�Oe����AG�z�w�s�j�w�5?�y:� �;E]���Q����S������E�W������}]#G�ͦc%���rw�h�����a�3�S��E�[,%mݟ��,|�fE�k�h	۵;	�z���S/�W���1���s���Q)�|,5y� �E������я<[j�p˯��oOܶ���q���EDAX7N�ن�]�tuR�qi%\R8�np{W�b�Z�"�oYA�D��,J���+��;�)�F>+�&��_��s�H�w��.�N�A�}��mF���������[�UX��D���w\g�q����L���ܜ���d␳�Z��Ā	c�qϟ���o�U}������x9w���dl�h�U��z096����/+b��������4�~�)�T9:�eOSe�Pz��v:��m*@`�����(���� /*�7�I�[)��D��C"��l���j�^�����S뭐V��3���<X�xO�I�I ���k�E�֡S{���6��;�*8�?PG�>>-°��1O8�s�Ō�lG�w�XJ�.���$�I����m`US�E��M��i�@u�o]j̰>-�'����&mMu�?�VF*�գ���黺�o�s��Z����,G��2k��B�t�t����V���؝:y;���:�nd��P	%��Q������V��~;&� ���FI�����!�` �Be�[Ԕ�h�U��q��6PeF��!L���A��S7gf�H��x���?�j܈���]����_�/#wWz�t=�5]82��>n��?���L7L�ֱT�(O�]1�
/�ᦳ	��x��Y�!yV�Y/
p1�[fs����>}���s\���g���	���p/�_���*��F�AI��D��d5DְJR����:�8�Mw���/����*���e8��4��]:�1T�(�ʿ ��1�Qȡgp+F[�"��,��b� �+(�8����#ݶ�_-�e�'�j��qRE2|k��?��F���<*�j�M7�+�����z/�����NO=
1�?Y��qf�H�2��i�lRca?')�t76�\�ls���Oυ��Ѯ��4���͏)T�..z�H����W��".k����|�RSdr+ǘ���sQ�$G�B}Xtr8[#+���!Q1վc�bbk��ʫ���ӅsNg��������.�2���w�*�K�(�*�W���_��d�RF��by̵S���VX�Ge~�<|�]�xe��E2�C{�'s2�#��@���S���ja���ԑÉ��J;�?���w��g'χ�Y�ֲ���g�c�f�0Q�3�������E�V���
,q	�% ��H\;MK�:����N�|�n��D۱��;̡A[\pbU��c�]	��z����R���ޓײ�"&��K�=��g���I�4.F���$D'�</m8�k�t�i��9?��p���P6��6���%����D���f����z��֌�Q��]"Έ�ݵ/���&[���ߚF�nG5���sd�ь��z`���՜0m�E�֍?ht(Tj|�b�6�d�y������2���G݊����d��L2���?1:�#�S�k�df��m2ۛ,�#C��>�f���[i�fO�m���@�>����>���B�{�b����U}߅�E>@[.�B�Ib3��:q��'��a�fb~xjV�Z��\�T<�ΐ��a��Zl?�2O�����'�-��r��{2���>T��>|�?�¹�q6}���|. Q��P.Hn&��!�輵��f/ަ&�2P�����k��ri�ގW�D���0s+sbSr�ϔLG�O�J�8A�Q2K ~gɡr�Vۼ�	��t)�����A�j$~��#w E���{�aX;�QZ�Aڀj"��?I����Q
�Ԍ�^�hi�;��Q?M���ͪ�^iڎ�6꾝�ѤΪ4r���ic�HY�:����������x&��\�ˠ��{��z.'d��묛�f��lZ6rQ���^:�(0�O�H�	Ӻ񷽦A�$�Ug�	���KWm��`vx���z�	7x�N�}besƘ���:��M�2T�0����k�7SB���e��]$�ƶG�Ƞ2M�dR7p۟�	�G�u|TK��e�ں]�L�2�
HNSp�ۈ���+���]�U���4�tm\�DO�E�;{��@3�B<��U[7�G١�E��nTj�Tk:[g�v0Q10�jO��t΁ɼ�V82�V��O�9rk��5/PN�6�/y�N�'�*1՚�������r��Q��ɡ��e���|�֫`y���uʵ�@�T,���<�@Nt�9,��K�"{1Lrhv����h6K�.�0�Mrdq�)�p$�M2G���f�>e�Rk��/D6���Mʱ�ǟ��:�%���B���I�4�)��gQ�Ć�B'���ozKН?
P�(�_�6��Sg�L�g)=�e<�����9u�ΰSK������<������v�z2N��"�>�~���`+��5�7�ă��">J��a�#KȈ�SN�`�����1G�8���"�ƫ�Ġ�x��J���ѷ���D:�K�n7��T?먛͏r9_���b w�w5��Y��Z	�*�/�=�7._�F}��Q��]#��@��+B�d���T�������Q(�oC������K�/�柕n��Ҟ�׹����r�eS�?E�{��VH�JY�>�k��O��#��O!�ՙ�Q'���W�������tc	-�� }nz�2�9Z�����Y�Q�k��\��A���c�n8֡*������ק\��mv�r����R�X����y�_۶��Xt3��e�5i��>[B�8g���=��$���:&�s�y������>Rf�q>n׺���v4鹜�qry�=?w��n3����C���_A��?���? Q�ɪ�6a�;��j`�Ϲ���i���~3m�wb %��:�L�L���
�}��A��1�����K�C`9�O��o�@7�����=
o7��a� _P)��\���r xܿ Q"�$��>n��Sm�I��U_rf�8���{^�IJ�G繜��9�C�t-�$҅��b����W��A)5����(�!Q��?T�2��^<���#�D���=Sʻ9��m
U������K��f�S�dO̎^x>bKA&��X��O��b��`D�@G�M����{�FɌ�L? ���7,�a��6Cg�A���(Ec֍w',k�՟�,;��Wl����[tW+ �O���3љ�w���U��F���)]�]�8<��&��/���@e7�I�����Z�Zk{��v6�E���q��|�h�h����ģ��U2 �MI�:XE'�+����_�)
��aASi1�;�K+K�sy��g0�L��6ѫ�����3;h,�j>��D��<E�{�UD����q�4&�� ��l�}<���#�&q/��>ř���P
�ܩ�'Ğ�I�+6@�W[b|�FR������Z�>h��q�g�񼯇�ߝ�����b��Ɯ�^uݔ�/����g�Yb�%E^���:�R�-J��
X���Rn}��`���oC��9��ʧlE���d��K�O}��6Q�r\�9�7�+��P��포�B�ܯ���N�X��	����l�G���P(����l�J�����!�l9���H���*�\>{k�q��H��}AK��"��r+��?�Ky1������W���+XAbDc�f�#���/��J�[�bu��y�G1i�J)���
�yε7�wВL��2�����֤H���Z\Pbm�ë��-�5n��+��U)��-��6'�㐸T�Z�M�]Ƙ�_+��n|�a_��V%���6W�x!�n�*B��J��g,l��Ѡ)�k}�wCM�Cdq���Й�1�w�\|���$E��џ>9��/:8r#7P�ę�{v��f+'.���1H<��'���2g#֖�R���.��J�M�yf��>�DaASN�k�`80����L4����c���b��R�(-o�p_� ~ۙ�hL�+�g��S`������E߾�c���Im�vL(�`��{���81�N4��0"�lJp]�.!���l[��T:mE��M0`�5�\�&��mY�f��������ʡ�7�L�ۣH�:9#6��?�X"p����r������DG�cR��Vdis$��]�&*B��N�ɨ����h��K��ą�i��K��ˏ�5K��!d�e��;���=�p	Y׬UZ:�����Z �Ҧx�ꭅ8c��:#V� ��eA�y����W�k��A�;���F��'@ܦW�Jؗ�u��O&B�:��t00R?KA��6�j������!x�u���d�	�Έ�%c��d���Ʉa�~�4gjB>$J^+�x�'?H����%�C��A�ߕ��Lx���W=�_Ģ������!��\�G)"���s�T�s�����2,���PH�5$��)��4e�?����R�.W�q�j૗�~�]q�?�;B�|_��῜�}h���R�3b�̺A�|�e�+�4@�Z-��bD]b�I�������p��E�a�%�v���QM_�@�]�7���1�B����QN/�����D�.EZ��X�X^�!8\,x���|��S�<� h�G��Y+j�����|��������3�� �
�Ɗco�(f�����`K������"����l�M	�2���)��'�=�&��Jԓ#bC^*&oO �>�W��X��\��U�k?��Ά��Lř�������K]&�9R-С�&!��_���	��#�L��s��b�����lCM���%��Fd%�v,���nT+*��4{	���W#N0�>�'ę�PQzK��|gTS�ҿ�r<�*�(��4!��t� ]��@h���j����J(J=�H�R��{'t�#�����?�k�_�e��v���<�L��<��|M֡�XV�����<A��6��|�D�U���i��iH��[����-�3H����ne\��/E\�e$����?��_��}|U��v6l�VH`�5�ז1�Ӧ�ݒ�j��6�QB|�� � L.�,S#��Q�v`w!�ZI��5��U4=�&���c��J�~$k���Ti���@K���~��O�{e��sR�-��(���-�$Gzk������^�iO�;�)��DR\i]��`f���,EB��'��g�=�Uh�����V��SQ9����y�X��@,�iD: �$p�����*0E�����j�(��h0oq�2Ъ�9�����qcrw6��9�L7�&�9\���]�������(# 侽Z׫FI��9�����7?�z֏fx�֝ �0��y �����)v-np�?�yGJ�i̒�=���`���!1a7X�F�í��*���>v�'$Bs�� �����$F���-/z�THl+���ϭ�T�N�@��&�\b�-����_6G�D���=>���)�5u�_9�#>d���0A���(�/�^���j���y[�%pH��y�Y�GR� B�{�,?V��3�C��X׼�P�r c�q8ޝ������(kJ����i��VHI������hw�9�Mb�>��l�jN�Cg[�`���$��\�J�3[����D)�!�ͳ��u�����fq���1+q����8�EN$>��<�ڞ� �u��{L�_=�-G��G�F�J��iih ��7��w�
ĥ��6K���~��Y-���ě�3,1|�w��$��*qI��;�&[��j(��H�y�9S$i�S��� w7P�Ա2��&'�����}�ei�q���w�W��{Vlڃ��Hb�z��]<r�D��H����; z]�����v�>L�%:f�6�`�kޕd=1l3U�����F���9P��Ʌ��(>G�ˉ�_��+6�"*�d.S�{Z�c?��_!�,x�绶��=�hH�bJ�I��/b�����5brʯ_��R�_AN*��Ai9ֹ���x���V�ON�;������~
��l�_��=�{�׊�J/c̸�[���Q�@Y���v�(m�ܴ�RI&<|3u�2�;c?Ѝ�Ş<��~>lU����Á٣"^�Ie�9�
lC������P�#L���*�s���O�^�-}�D��H�D��S�fyhM��v#�͙��e[���h6�j�N@(�e?�?���3�;���wF1�40_\sV�joe���׉ ���}��9�{���Y�~��I^�2���/��|+�����j����ҙ��w^�1ryO���b�]Ӵb~{�|�yƺ��&�l͹����.�q����6�`<�A,����B7�$�4�1DV�H�S[�)��(}M����f_.sq���Щ�K�6���;*�]ju�'�������0&ѓ6�g��?��ҵ֍I��k���b���j��9H�0��?�}*
#�Easn&��E�'k�m��vJ�/��yu���R-L|��%JK��h�'�3L�j��:����'�P�ӧ)�p��i��ީ�%o}2�t�|>e���:h�8u�e�O��בݩ�W%~��_ݵ}gl�9�@���,V�wVP�ӌ��B���Qߟ�sA�	�3V
�}T؋L�}��H���V�5g��5i��Իb��\D�<!�ǌ�.����Q��n�k�>�_>�u+ɢ���&z�����׾4�Go�p�S��+`��j{v�FoEx�
J���a���1��ԊL���!hk���m��޼���g�e��Q����齻���%d��^�	zb��fb���_�G�s>p
�$����ck��ɬm��ú
WV��
�&G��"2O�T1~JOfW5M��ΊSc*@O��7����bؓl�12<Ŏ�0����!O%|�Q3���7ν]N~�4r�CԄ
�(���<�
��!ZI�7����E�s
�Д�ɮ/�5Cc����<DAN�:��U$���B^��	�����9ܚ�����[�1!]�A5˝�-�Ԫ���!���<)�j��2�K9�q][��ػ�+�K>s��ïK�C!G��.��db�@��#+A<֨�[������s8l�,7|��p�͛�:���񮢼��Rc;�Q g-VO���	g��ᚾl@�ȎSg�N���qP����`�-�U2(��Bxn���^�ZB���w=�I�t����8(��F�Galu�Y��\�҅ ��bP�E.��3���?.[Ⱦ��h�n��E(��6�{�U3��V���:F���U���L^���;�����>"�xD$�݈�Z�gD����n�l�p[:J����у�^���*E徕�//:s�;HK��&���ļ���yy������y�m�/��Χ�PC[Wb�猯u������H�#�g�T�y�E�Y�ce��<>W��:��5�Y�қ�"_	�����g����n����8�n�nK󕼛��*x��Ss۝ �~n!Bz�מ�6��-f[����[^�s�� eM��MǼ:��r=��@��F��s�~���j2廬�M�7��E�|&x]]'V^�����`v�>�B���I���V)�����2���I6f�l4=g��7*4a�� �>*~⺼�H�pIM6�-iFm3�����]0[��).pA�u_GAAM��P&©�T||�kH-4=�:NE��8�H
296����Z=~����^7-��u�~>����m�ys[�� ��|2���E��+O��kq㥵����b�N�V_�&�˷�r�˴S֬��ļ��ng�����WE=�\�rݼ���6�ƻX���=�|��#���K�Yd~S���{[fl��AȤi��;4��� ���Ҋ�.����Y��-�f!�e�z��������Dw��+�V�6!�>�|��xW�ڞ���B�aޜ�a=&fEҾ%�w��H�N\�
q)�s83��U���<ٵz&���:�*&C� ��I��T���wW��t8"$DY69|+M��w�辯���?7q���cZB� �ķ���F	���᧪������x�EQ]ѓMz��U)爛t�B�6N?A�ֽL�`C���w�_-��EP�3E��N�]M�H�q"D����HI{��3w�@m���jF�$�6�ZJ �B�yx��-�Vi]�O�<S�~�k��]�.�I�+���e�_v�����z��f�Q&��{(뉡p�+�s�X�����H��B����j�"5��|Zk��$�=����+=��?`4l�k��"����=3Qx4�ܘ;��Fn&]f�V���Q/D��z~գl�S]ct��ڠ~:�h�s�l�ב�Mzѵ��W<HSUiW���.��aH��O&�0U߸qRk�SM&�i-�yxńY6��˜O�5!�Y���<�(����E-��=�~��ˡ�j��a�5�����ƩU ����U�:C}vaf�Z����U�e����(�TWTjm�*���"
j]kڐ#B�Ć�V3k�^��U��wbv[�R���UҦ���b^!܄�xL)7=��<Q`!��9�9���g���&��ز���u����(l~�I��Oj:�*q�-C�x��[����d�ƅ/o�sh�
��m�C��^*���yB�b�ʑ��ؼ�`��B�\���?*��8�o�:�vU���gy�)����x"ڋ!Mc$���.��V����<�v2�mF	p�9�'�f����э,�vj
W�����5�6*�����ٻ^D�ϢۣD���&S�Pz�)vz�dy==�����2�a�5����M�:�������p���Xt6N�3G�0������c�>!�UI)z�X�~��YNs!���86�]����$UtK��3���*������6�\���+`�xU3�UQ��#=->FnU͒i�I��z�c&�҂�i=	�[�����i�ڿO�f]Ii=K1�[�D�A2b���S�]���"��
f��a�����Fs&��E�9�/�!��]&�����d�J�=����V�����>G������r1P�E�x�A��za�����(f���0*�F0^��c������l�sE�Rm�������Z�ΈL� 0�e���!�*�>�&�N�BG3#߉:���F�4�ÖP>a;�L~iɔ��u�lhk�UtWN]jdcFsT�̚e��`٧
�i��}�Hk'�'�v�)�0o��=���ꅽ� �; �5��9A%�-�3��C��!��OMY���)��՘�oÄ'M1d���j�>0�vǡ�FV����'JJ�7^�d�K��Y��Ĳ�d~Ď���t��w)����e{�l�=���w��,D�N]��V�A����Co&~2�����d�%��r%]�9�_A��RZd�yv�L�w�|Z�?��u��f�BP"(�Tm�6yS�s�,�t�!f�� �^���e.�5�ɰ�/B6MW�>#N�ڟϷ�Q��+�MNoǐ�<�p���;w)9�T��%�y�%�w�`j8c����Y�SȔI;�ku���ܪdh��'!�l�L{���F�:�<������4\��v��E,�;�݅�Cx�./�)��.�����iu�����i-6��j_�;n��g��_>re�oJX�K�27Z=�u����7m��ڊrǂ2[��:�p����id���@�D.)���o0��ZX��q� l�bTJxs5�FN�1D~;ʜ`��j_'!n��y����XH����2��qO�к;VD9��]{zr��z����T�:9����t��M�a�:����r&�I&����Q�����up�r�o̠;�x�茪r͢}���3t& �縶��Eܕ .RW�\j7#no�\a��v��E�v�yr,�˒.8��*_?ɬ��厏zsಭE�؛�ͳ���<\D�f"�<$~z��N���y��_��Ȅ��/'�
�X�ŝ��G���Ε�B7zu�����q���� ���AG=��`ŪƟN���Z}з&b�ѕ���[ZY�4� �i��Ui7��b��SB����\���O7��6�%JZܲ`�������ycD^X�90퓺%��3��@u{=4��*#3mְ>����Gh����)�Kq�f���ex��k@��r�5�2�~���"�eI���L�E	d�|#E�vee��&�����:aj�s��[q[����S^U���B�bEN�V4�v�a��\T]�3�L�߈/�jh4�H�Zv`�X�G����2�q�-��b���<����c�l��:.���L�h��N���K�x�!��2-�:P�)�$r�ʺ�)*q	�mu��XM@n0�2M��ݍK�)�\���f��y��{uP)�� +�{�d(�q�n�Y�BT�c�.�	��2<���lz�-P�}�Y�
,�P�p�j��q����	BH;�P�N_o+w��2��(�0`�d'�9�**���f�9�U�I0���@N9r��
�������7�l!6aT�9����Bp�ԟ�
@q�|�i�L�OL1Z����H��ۢ�r��3{���]��ʖƬ#��g&�DA�V+�"��{��1�	o�(_����T7����(��#���L�c����Π�O����:��hs�\+�jZS���u�����?9d/F��<�j��h���D��U�_kDܪ�v���L(E�o���5���֐�<����\�0��k_�ݔ~�o�df��|c*��&Ҵ/�t��'����+��9��:�'�eEy���.`���x;�F���0N�wI���1RW�c�W4,����	R����kgZ����D*ՙ��fɻ��c��GX:�^�͹���}BT:v���@Q��Z	��gdϣ�q�[�2����\��+�}���W�~�<j�*��N�$�@ԑo'y�!X�l�m��Ê�q�@2�5�"�����+\�E�9"�� _�#y�N�F&C��Gt}orѰ���D-�r���l��-���<����'=�P�eq���>�K\���(�S|A�7D����"$5h\�h�z>�N��?��S���ʂ��������^�$,K�Nȹ <��/Y�<˥�4r_tg��(&���I�0qd���"���i�
��g�{"�b�o���C.޷�~d��$��3����}`MG{ &�E�25����Ĉԭ��M l�����	Z�g��.ўrd�r�Ϩ�Ѻ�gg�ý#-�M����w<:�}��Q-�b\?���w�K���d��m�R��YJk(��e6��k����KxH܎^8{���3�[�i8��%×Ff꙲T"��x޺f��M���3@���$�����0h2]�G��+�#���a�v���I��Yқ���D�q��!S}'{x�ی��th�-*�ś�w����g��@�y��V��BL�e����.B ����V��"x��˜��] �+*'�a��M���*�����#���s�c�A���Ğ�~u���Y�ۼ�1��"��Q�ǂ*0�`�H6��%� ��𲎔�N�����?��ap���)��P�}��	����|-u�� ue�%��I1=j:8�~v���[�~d�T�*槣�c�EPO���X�L�n$�*4Z��o쳎o?
Q�T��|HA���ˍ�oϥ~�g�;��2q/�������\�_Ey�������P8�s�bɻ�ĝ�)�0&B(�E�z�ü+��-/?"#�E���[5a��%�}ZZ+ e"Doq�g���'Rm�U��*�����U�Gb$X	� �>�͔S;Y�`$��U祿��r <A�r2��u������#��̇9��W{���"�K`.Xfa[�U'ٜ��R��bh<��{���
R���*�* �L?>]��L:�Oy���Ot�^►1��b&(��*=G�6����2^~��s�VM������K�1�X�����|��0X��9�Ogz��@!ޜ�0IJ������M���u�}['h��ow&�_�hO�)��F�_�d��
r|k���O8ߪ����CF[�E�	�J���!��ʕ��Ǝ�/ɽ�������ukך�i���b,� ղ�pkB����?���x�tu�DЭW�PH��1'������S�R�$xxU(O|W�Ş��Db#i�����<���^,���Bo�"���HuA�2���#�i��F-YC�!���K}�.+A��P&¦�����)!'�ȡ>s�'9��ݥ�jNsO��QcC��5�eI�pO�◱�6���Q���`��	�rLaM���m�Ԁ��%��lw��Z��c)ϕ���y
L��h.7yz��Q*ɍ��S��Q��l�}�XIe��Y���ɩM ��i�e%�4�y�_���	r��LE��E��!j0���ɲ��)��S������`׆�Ǳ2ޥ������d�,��[��.�窘�J��7�߽���N#eRǢ��ɳ�8��>���	z�q0@}����j]��l�t>�)!_(VX	ݺv��V�4E[�N������3 �������$_�.��"j�����Jd6^��&�~�I���I8�H@$GT�&�bˆ�Id̲(6]����3m�[�,(,I4a������DT�k�?�\J���=��(�K%�:Y�H3�u2r}��h�׼
Q��u��m� �82"����%��L���%M�����Ċ8T��Ha}���[U�dX�>.�6+��'��tN�ʖO�ٰ�4��ƹ�NJsEa��/��~&��W�������L���zD�!�-i��1?�c7o�aR���:�SGg���pY��C+߰N��4���m����CZ'��N�I܏�_��4�i�C�"�a��Ä�$��Оqn���Yg�m��Z�̺�����'�{�V�+��f���{.M�7ʷ�G���135}^+��B�z��o��ڠ�Bo2g{�>jwb$��Q'�̐��p �7j��PX���[p��r�Aw�5e��M��W'���������b�1�n)^[F7��x ��:�����/iڰ������k�o����A-�\��Ǳ��؋�;�ͷ�pK��z/{wk�N!���V��Ҹ��u)i�x!m�������A_�F!s����?�?���_����G�/9S���ҭ'���8�������N���H1���?\��7�s?�$��_a�}T�����\b�l�255��7f��
`y^�N~��g#�m��r��|�;]mdĠ��myy�����NNN+�!��1��k+�h�����Pt��eT5���P�/���b���/��?�1m���������_�/���b���/���O���˿p��RCE[9�����PK   ��dX`$} [ /   images/a8bb870d-02b9-45f0-bd60-404fdaa8f6ff.png켉;��?\_ϣzR�'B�OE"b,-�����f�v��Rc�Z�P#$��R�l��3�c�Ⱦ������{����}_׹|���9���������u��;v�Ӿ
7ܱco	�{77��'���������O��X�y���[�;D>��wV;�0�Bk�D�ۡ1V^�;0�YG7g�����Yw/�D���;��І_�����D����,.����? ��?v�@ў=r���>?Ot�8���g�8�Ko��ve{��;��M��g�d��&kܖD<Йpo����k,ѧގH����@5F�G|�X��9�@�j`S.�'��[��ؿ���\�m�݇m�h��Jx۵9w���{�D�c���W��%\[����vn}����ma��������Ƿ}>�cN{��!������	�#�{��.��26��������.��qDSx�v���61H�~���/ڈ���V��|~
t�Kk���!Q츨(��?q6��k>�4�r�K)�TnG� ���*�E�Op�@�]��\�;/˘a�y3D}?��J�������%�����ٌ�<�U�Rb�pT��f�%�\��$S��J�d<�T%6��#AZ���ǻC�zs��0���?Y����z����c�*�9���ޟ(8B}�Uv��K�!���W�DzS�ڿ�¹QFn���\-�-|�&L���X^�M֫�-�d=꼒��t�?�>,�����3�ah�1 Qf��qːY�����)J�	B|U��"����;h�5횇�p���7x��-���"ǵ0�Mø��3j�3��$���6RɟVS ���Y�|䟇e��&m���>.�E�{�.�Hd�Z`����)�E��w��4	����ۦ	h��;���b(��?���3�nԛijiY�7���[�f���ʢ[�M��-o`+��]�S���ḇ)�˨4�`s��ϐ�5��i=ΩX��\��0�żӸ����Kpx��J�e�ztW�J��erC})�� ��s�>��+Ȭ�?'�a_wu޿fg��0�*�{2�as����@ۈ̥/���pK��~p-j��uۖYo*�%H�Ab$rp|�,���6�FX�0��y=�M4n�G�'�s�_�e����>���x�d�k�������f��$�D�����=��_;#�z���c��$w�����O[�&�V�
��?�ݾ��|t���A��U���à�Ϫ^&��A��uص���qX"����
+u&��SJ�V4S8(�}�")�+��i���k�<j�~-�=w����1#��5�E[�ws<7:)e�wmt�U�#g��r�1�jB�{	*C��/Z�X�����V���E�i��Z.���E�pa�L�PS��<���w��C�Q�S޹��G���)!�*u�nˁ7,�o�n���b�:u�J�����f��A��J��'.f����O�-�g��8B��$�PI�7u���;����z�>{V����K|��Zy>A5c�
/g����1�Z)6T��|�/*��,����MD�8֒��9��++�����4�`z�Mک��e}����ќ��CYI���
�Z���ŤTe0-�FY�=8����E�A�]c�uc��^�/#��F�R��kqbi7�jԯW��U1m�/̏��bh�u-m��y���W>-�2�߇	M�H7ڈ�2{N����b%�뜈�M<�S$��r�Ot��e���K2ǯ*�|�í��������'��k�������:��a1�����J�����������&�#�&W�J�(�bUOx�J<v����.��rcqC#ĉ_�E��f|��%�h0L뻸�3a}��a�k��M���<^���~(���`'���"k�	=`��5�����^�o�EjB m��h*��ɡ�{_��'x������R���f�����Zm��f�4i�U^��AT]��!���Q�UZ/E����ÁD�J+��նܰʶL�%H~�;�g��ƢGF�L?�����ť}����ōϦ��?ʱ�c�����d���^������k�i���IL��@�dh27N(��ԿaUJcmm�O��y�w=,0OL�G
��;~|�*��Kc4��M�7n��`�c\�����g���Q���I��Jg|f���v��h���)�՚���mr�)N5ڤ0�e�X}���{Xm��_�ƺ�"��%�#ǚ�a:��$m��ŗa8�$����N�B�z`���|
��q�~���A����ӻ=jić�Q}{s��6[�
o�J�$���j}�~��P�p54�!�3���A���F}�©��S��C���q��9]�OPY�v��r�Y�0�gD�0��gLm*+�`����pS�lp�����I�2�rP	~!�̕ߔE�<F	n�g��a
L�)ݽn��}����B+	e�h�s �u�L�j���n�t<,�M6S������-�2_��+@�p4�Lʾx��^����p�U���q��ҁ�}!��Ya�� �Q� ��ʪ�S�oC������������l��Okx����m����V��S}<A�mH�\���E�ֿ-j0D�:�̼Lڸxh������e�T����Zl�\7�I��n~�b77�N5i?[�SlD���6��$�pJ)�>x�ܰ6�:�v��!�	��J�"fz)QÿbJ��@��N[��niI�jZ�N`!=>��#o-(�W��\�:Β���	�9�qyӒ-t��4��v4p+��a�7/yF�0�#�j�;#�@�_2���q�B�J�Be�p��?4��j��n*�����3_����j���*�~��v���7���m5�i�!�P�V������P7����;~�M~�2=W�q6RkP��*��Z�>r�&Xryk5,�6�qJ�ϖuԎD�z�K��򥹇�+|�XP������HY_�(�X�ԭC�Λ���B0�������c��f�M,;RP����vQ儅�&Z aa���7��F�r�=�Qu;�HN����a���6��2�\��,Iq�5ăj\���n�OPa��)_Ɏ^P?���Iл�CS�� ��n��M��f�F�AJ�Q�jhȢ���1?P(i!2��"Цx
�?��iAH���I�8���5�Y ��a�|�ƽ�O�:�5@;`2,�1.&�M�hh�_��ӿ>� ="	�I�#s��ʝ����������k[���ͮ����ɗ��Y��6(�_+Ps�zuW���k�y���H�'�v�����wN�z�7���5�5����ˬ˰I@�X��&˿G�(�4�0f%��O�#�e1���
G�3�w�8fU�Y�k�g�6��M��m4��'��L����*�G�F��|]��ߘ./�t8�:oYԾ_�`uRRleŋQec|2�=��W0����<&��"��t��I�؍�6>tk�����R�|�U���񧒣a֝�,�^���>_jo�͒��7�� ` :OiI����X�C��|�_>�$��$Ptl R/��л?=�;��g��*��5�
�UN�s(��w�*Ս��ΟU@����+��*G��)���Y�x��%vUލ�X�uS�"X�#'P�O��y�_�r6JB��7x�~b+�)⑰��&�G��[K���ק
f�<�'��N��y.R,�$bΧ��ʬ�o|�:�g`�v�
s�	 �wp��e���r6�Z<�	��34U�_/��2z:rl҉�F�ޗ0IAkv�̯a?�r�b�g@����i�	�j�N�N�?M���_��I�I�KD`Re����3�z���T�����H�@���
���i��G���������z"q���Hni��}�Z�G
�,��)[�=Vi*�W�Oc�*�j.����t.�V���,�t�a��
!7S������䕘�ƨ�5d��uX���y�]Tpd��LgA���`�:xgh Wm��n���g��kȹh������QX��+�I���a�kډg�z0���n-�Xډ��xOh���b��Sa�iz���s}�������l���8X�ZX�}u�<�mpT��监�w\p�Mi>��=R��I�R0��J"U�0,+ng��IT�FG���C��ɭi�i��%���r�9��\���
Ǧ�-<Ş���C}�~����f��|#@v%cBLS�� ��[P�����;� c��=���QS��_|ɓ"��A8��6H��X�^QH��t2�nn��װ��gp�V��Ν�<qh�J� O��FIH�T�<	6�`^-(X����v��V��>�����%�;K��Ò��t7w�DPn��[��ZF�[_�8�������H�\���ݘ��0�`ב x>�[�\�⸓�i���Q@#�C4���7Pk#x����F(	�/r��X�����ɽ���D�j�| ��k �z���c�$������yiܸzE",����h�C�����b�b���D*��.�������[]��\��]ӆӊ�{V�VN��0���5k�$��Ha~��s�ﬗ�ޘϐeW���r� 9}����f��i�vn�:T��in�R[kq��	�1i�|����ˤTN�O��U{u�!{A����w:���l�դ~LҒ��\�� }�!��|\�I��Y���$/�v���ԓ'O�񰱼��kK�Z7�H�W��$���G"�0B���]"Gg�ċ]�.X�;n��6R�{��Q�۬p����G�'��f��6�:�w-��@��>�)iii`m%�^$�\��Bx���I�ŉ�xE�������N����œ�h	�+�>�uJ��D�0�@�}�����]��}ݣ�k����%�A�5j�nq�oY�\��a��Z�8EE�q��u��E͚ C�TV���Y�S�҇'�I�,V$�2[�E:M�my�D&?7T�A#���;�� ����5E&���4����,�;�4�e��̦��
0��,2�v�|���ŕ(6,
��s0�E.�Ҡ�IX_'����9:1U1"[�ն5�;���_��R���u	�F;��uQA��������b��L�'�u�'^�����J�ƀ	se��?E럼!�>���r-�5E�]��h*���!��i�#4�ҟ%������YS����J$�=���'�L�Ȯ���SƏ�
��/.M>}��\��+nll��3�,�=<~�b}u�G�Z.}��0�}" �ɹU]vʹ&�����S�FK�<4���'�]�xXZ`�T��_4��sW�b�VE�2`�b�88{	�T�AS ��Q�����,�g�䔟ck�m��e���P�
m�.��|Gn�Cٰ���TTֈX_��"��'��"JӼ0�a�{25���6�Ȩ�_�2S�k�m4V�[[$c�� �[j�)�m��q���R�,�R��D.�.%{��b"��ݵc�M��_GiJv�j3`}Ȭ�s�T���ӮMz�wԏH�O���7�R�Jt���F"M4k^���b-��5�y�fk)?��Ł
y	��x�{:��V<�r��	�5�>�o�fH�T�H��^6i|{3�,�ɞ�CV����c�T�e�8a�c��d�>��Oi�.�9��=��d�Xt8ȫ	@��a����j��H����z�.`������!�Ҙ}��U�E�1�zfY$3��Ėё�Ƀq���#�'��@��I$��d�Lk�����`R<M	6�<R*�z�7��x���jM�iv�my�?���,�nJ{��Mk��|��0{�����4@�@M�8�������[/��Q_�~-�c�ӄ���OeB<�Y)�O��ǉ%��q�L$�)7�)�hm`��Hz�
�Z��#�/�g�zc�{=�B5k`Pky�ѡ i\߉8�t<��0 6|�G����s�X���E:�$8n//��Z�A��;�� $��Q�؊t�� �Y.�bk71��K��s$��#�s�A������W0����by���vS���.P�ό��~ rK�$RJ����C��e��\:�d��W-�r� $7��R��,��(.���re4�:.N�g��g� ΍��{����!޾�99��($f�Xl?j�Z�LR�t�m5�2��gk�ɗ?g��DJ�1 �Km�ȅ��j=.
�C�$�Q���z��m�C��b�a���D���T��)9�ڇ���Aޢȩ���� �b��B�s�髬G#>��ֽb-��1_�)fw��"�G���K7�< 5݊�-��6K/A���.�*�kTK2t�������K��W��Q^�@D;�L744d�dך���� {�B�$RH]�5���Q�cw�k1wP/��}̦l��Y7��� �!���.wAaasd��~�܉���5���Z�p19܄�������ȟ���Q�xc�����Ea�A!����-��3��r:2�}:B�O�p�qz� `\�Gр���TTk�Q|�N���E�e��j��}�#x���� =s�q�R2���	��!��w�:����#�y���Km��	;�/�a e�l��J�-�6[w̖�#�.�H�Bb̫^��gO��Y�PX�o����<�dl�������igC��` ���6�Y���"��{�7dz�K�GtN�ⰦR �w�R.�-<68s+fC��Bv����Q(@��_�re����}�kG{-^#μ�����9�Ug��y��I����B�����6���.@}��R�J����&��L��T�$�Te3o?����H�c�7�ˎ�v��թ���ї��кHd�FM(�� N:���_T΁���l_~�(�8�\KW"��H���D����l{:&S��pǾY�8���xq�}�P ��i�E1Щw���,��
��O�H�D��k1��V�`JN[�ً?�t�9T B�.�4=̃u�e~�G��u��	��'�Q�F�4�h�$�5��H�q���	��%�Z��g���u	V$�o�i�ȶ������ɔm`�D�����)��Пѕm���H���t2 �q����r�N��K�������=�BI�E�"�Ͳ�ȨPU�yՠ�i$RN��	@���j��h�yS9��~�b-�x��}���Z�J�ċ�ۦ��K��/N�3M/_��,�,X��',�dh�͏�}���[�@m���\�a�Sah�����{q���ĜQ���]��+�	 ��H��E����H+P��L|d$`��keJ��P�F�s�`ˇ�-��gP��t����\���R�>d:�9U ���Y����ר�N*�������A3���� _Aw+��0�FE�Ww1�r-���)է��2�E�M�/Lrn/�I� D�~���d�"+�ާ_���Қ�w��
A+��i�wI4Bd*��e�?^01���!�B?���P���X�B�� \����#�&��4qh�������,Yy��/qQ����k#o���[l��=�c������zY@��W��=b��~��b�`�L���'���v*\��C,X��-$�!!�/����?��K�wp� �R�kj"l����-ҹ7�f�A�(�%�#���6	_^��5��f�k��ɴ��s]�	�%�_�;��Ҍ�� �1��:s!�Ν;άe&Y�e��L����$����������9'b|���+�}�)	��ሺ8T��rnn��d�
<��)�e�h��|�	��G�}c?����]���Z�<��ZZ����\)5;��\��K�%$�4�����\���i�(`� �ce���0\)�I� ����?�gs�Y/��T?��j�F+EQn�۵�Ҏ�E��ac�g�Y#��b���Zkw�_/]��*
h���S� l�Dأ�<v��Nv`Kd�_W%��y���f�d?c�\]YI� #�^	����-K�av��K�B��p��-�_������-X�/Tm	� �)`�|66�&^@�����,T����G��2/���{�����ۥ3��W������Ȋ��[$�w�#s:���Z٨(�7�P"��w�~�n���A]�BY��sB��F��럺%{�h�P���p!��!��v�����8EY��nd[�.�
�z�4`���HDa���fw��e�L�* :�L5�f/���"2�� M��H�o@��D�,=�Ӫ���\���*y+u�p�v�N���CM�q%*���v�E~��M:�"A�b�����@� Ѹ����N�� Ye���"���^
������VL��� ��`K؎�a�K%kNo-���/�����Rs�~�o�v�����3-R�}����0��#��r�i���e�i$��k8����=;<����خ��W+V��>Cd�O�>���\i%ӵ��h��Adk�b>zע���"(��5��T�u��d�f�)~}F4C�#��)"���FsY+$Ҽ˩Э����Ъ�����e5��A�U��'�u�VCj�8��$���[99h U�J�A�,3��0���Z�M��m9�\K�L�]e ��]M7a�?��(J�c<`w�s��T+O�s�^XMi��g��?�S���-��~du��V�$�@�[�9 B�������^��%���H΄���<o��֒,+���~���J�L�U�ݻT,��+���؞��G*����Yv�]ߡ��ɲ�~�tځ���[s��5�j�	73�{�-i�(���P>�[�KMS_K?ӴWѥ�k��矠!��I�Ǳ�7J��8me:���pv
A!��]��2�	M--��C�nB�3K�>/Sai@��=מB��J��I$I�]����9�I�6qi�a��m\�_y]X*yrxC�?�T�$0ӄ��O%m���fAC����G�@Vo�a��gO6�e�Т7�8S)j�|��0��,>�~ z�c��r��k���ɰG�@UHA�b�=���OF�2��=��H7&�Z�"2�$�q�]� �G@0MJ7���]<~�7�teF��P��d.C�Lߘd������+��L����w%X��`�tg���}����L� �n��y��
�
�5���WVn�/����tӗ0O6S�O��9r���w�O���u����A~�2X�j�Gi��Z�(o��7_���D�����w��H��(�$���`��	�6U%�lR��[��T�;�k��-P盇!S��Hm��Y�W�1k�?�M��n�
ǁ}9�6�q)���+MM��2�;õ�y:
v��7� _q�k�'}V�c��,�kV:���]�]�P�_ld��ڽ�5�*6\�d�A�ö�(�"LL��9�F���-�Λ�(�f4�F`�e��^�Q:v/��trm�Y��`�	ɓ���d?���x��S���ט874	�5�]Q�i	��N�A-�R��*����t1a�7]Ry���yo��b�V����Q�1m���i��"B��A��ݾg�u�Ud��	�����pDc���!@�Hn^��_$��<��&��p"��)��(�����5VGZ�I�����A
}gT'����F��11��ͧk�m�N�׫F��4��I`
(&�0?X�Y��`-F�7���?3��n��(���< %�X�Qp�6���mM
܎�D�c�(lCo�}&���9c�ȍĆ�0�Ȩ�='%�eO�{����wf�z��y���î�j�F��&o��x�Z�zMP�6��'��[�w�t�(�BB@2��:�A0�v>;4)�8�H�I�8K�Ȉ�Ol�Ě���:��P�+��Z;$r�K�y��{����8l�6z���cn�~�{5+��`��'`���yo�	\��;\ó�"|��M���sd\�%d�;��~=�L{6eᰋ�x�4��,�����k�DH"�<iR�!�7Nb��;�x�5�s����a��Du��Y�Y&�1d���v����1ZE^��6�;���*��7�}�)v� �?�K1�yw��8gr������n��b_�֠���V��!�{1�ʊ��X��M~0�&˞� �S�;^��t
:O�{	�c�nƍå�y��/qLm< �� D��ôgh;m���V�����g����Z�"���v�ç�eN��D�n�8/�T�/��]K�/���x*� q�C��&:")����!�M�@y}?������G�ث{]�c���H�l�����ɵ������ɈL�)�t�C�+c���.5j��|z\)`���OC������c���+��C��?J�)ʌ�@���]�3�UΓ���o/�O���%���l�E�Ѷp)�,�ɜ��|�_W���'cX�YD�;eG~��Ću�0����0YѺK�s����Ǖ��MesU�QzD\�B��o����	}��1`�;���ՀCBҬw�����U(�ΐڣ�����?��Wǩ�Wkf�[<���C""��@���VN���h�����= ID`x��W�6�8c��{��Բ�;�7�=����LV��&y9��҉
D��YUl�����h~f�jg���~�sU�n�5� "{�a$67Ț�����uU ���7�E��;o'�̹����_}x������e�D�_2G��S���y�÷�[��>����`��n����rN��
w9C�}��9(vH�t�,��V�>NPX*Y� 	��W����XZ=t8�*\=���y�4�G�fu���e� ���5*�Z�Y�tl#\��5d�+Q��/����V��l�`ĸ�{�7lt]I��RU�f~�nտ<��0!Q��<��x�NF��� �ͱW����]�=��k5-������;����'��|L�(�m��p��j�^'������/���Z5Q Y�����=��1�/ꞃ�����{/���s�Ĭ���VDs-������{OZ� �T �vV���2��o�C���6.jj����%�t������XJ)�	�q����?�4����2�$iv�x���X�FxxlN|;M����������F2f�� \E�A���j�-�DI-�^�B��A�����	h*�Y�lx��A��	]�d7����g|�8Ju��rƩ{K"f[���TF���'	�HƓ Ti"�D �,�##���,|���ԛoO����و7-D��&�U���l`�'tt�y��\��A�*�$��]{5�� ���5h��	�"u����"?[��: !D���3�����@�Y)JhU2Su��� J"YHH�g�뷙^��Ei�U\u�F��B�>��ް��F��������j�1P�ғ�ّ�@/ʾ�g�b��>���bN<-
�����e;���S��Mi�,P��8�ͧ��n��ڮ��"Z�IxC�2.;���F��s�Sp�ǹ�i�k��'���y	�3��X�C���W�
���h��3��g��B���s��'슨Eٝ��g�W�T��ˉ"��~���L�,l		���#Z��uIS�Ep�O�������WeP��֤�����F�C�ܬՙ�]*�����e;�껡|G��w�%�S�w�Ş��pǏ��*�1�S�U;���(�����*HT�W5��+h��:�/u��D �M�[���T.A������pϭ�/n��{0(i+zx�>�[�������$��u3�}�q�XT�k4��M}�(�������4{GJ�X���a~o�n�ĎE�3�-�8Ne�j�*�_mg����>p���>(��L3|x-��f`����p!p��+'���N��x�{�M�$�=�~JC��^��4x�l'�/Ϧ^�eԎ���+(1��YQsγ�9�d 9v�*Ψ�A�n�P���8!�1���H����o�P{"�3����<э����޹�7-
a�^����\�;��DJ����E�B�G����;O
��w��FJ,,�~pdR�x�=O�����[� A�T�M�NlB�4e<�S���k�y0�#��+=3F ��)}���Ϛ�a)sNm_�lڑ`�Z�x�-`�/9� �[��l"׫���d��L�Լ��L�U�#�^��5��L��J9��
h'�iij�Ĺݣ$���q��tT���hJ�͡�n�.��ەq�5�Du���Qʭ����ak)�b�
5�y������*�5ۿ�����$Q�c0�P�M���^��.9�r^�����h7DLL,�����=�U�
E)?�i(!g�+p�UF:�oZ���Zp	����7�JˍRhk,T2��D	�mkk� ��oy���������E�c}���aC�d�&���aZ�q1%Эzgؗ���.+�ܩޙ2�{|�����}+Ľ�� Ǯz��q�;`��������zRB%���R�ͯ�r�=���9R�- �^a�o~�j��)͠E&F�/�f>�%�> N܅�_c4��B�"�cajg����-��ph�FʜR�_8�֋��+�:���ޝ�+��FY���qnY|�����=�V�)���;ĳ��+�����_�H/;�,	�￧4����ؿ���D�T�+n�=�W+���F
����=?�d�S<ـ�Fuv�"������Hq@�>g&��^o�Z&�/?���f�%'�Uٱ�e7TԚx?Kb;�+,�j'
����p=��eN�d<�w �S�E���$�Tn��6���J� {R.��Cvˢ�T��=��JXJ�J)u�u*����؛7@ϔ���LKB�J4�Ji?�.'���<`��-�S:j�Q��;NL�ƹ	W��s��WM)eyEC���3��W#y�t�cz�*x��6߃=��Cc�MD���5W�?���8[J�*�@K�˾���0C��Vh�x^��[�s�����p�	"��D�I���K�Q!�s��P6o�w[����3��)./�ͩI�~��cH[ʕ+V	R�>�xjݩ͊��
���dq������;����3t����d���v���8U�ک>�/���`����,�~�?�}������P�	 e$6lo�o	��io��K��H* e&d8R��f#�l�׺d5yn֙�߿��j����U'
���DW6,����SKU�m�'�4��U�`jF{�٬�#ǮJŶZ2KT�(A���r_��KB������o<������V�y$�-�FE@�.<�-��撐���r�Ox��aWZ��&��Gt��L���!U{��t�h����P p��ȡp���_S���#�<��X��e�ƩC�Cf���N8���ܕ3�y����o����a(<<�`5�1������j��>�A��j.�[U?�Ҫ���	��[�[���
��`4
���$�Vl�[4��j�v�ߊ����7m	�D�v�(K	�̻��l�-m��y��R��4)��)�Ӫ4��]�~FW��[7�1��N�8V/�=���Fr���EwP0L�R��R���t?����?�9�Հ��xR�D9�;6"��d̼Z�O�F�&t��q�|�ʵ����Q����`�y�d�ܨ<�+�=�պ����f����.��~ԭ�(4�������z0^�>C�Y�pB��� �����!έ�H�1�{/��h�2+�WX��*
'߃��P���_��}C�Ȉe	�爝 K�ɕ��j�H��!�����/w��l=�˸��&	X��
�f�>�>��-�Ů���حP������|�G[�� ��t�D����է�aw�} E/��)o�X�н���p�9$�%|��䩃BH&�s�#��D�=\�
�5�6=o����Ha��!H{�m���'T4�6� �.�DJ�qq����(w��N��Ib!�H}���W��[��� ���e �}���[S;�b!`���?{t�PbXFa��w�2䡅~-�52�v�l���������A]�ȳ���6l���� J��yL�90��5B0G˽v��DGGFbOaOb�+d������� D��ֽwd|��n�����`2���e��8�!�����T\N<��BZRxg�q��x>K�)_�z�P��ȼ��΋Ld��S���q�w���� ��~������U7f�Ǆ��X�{��Ndz�*|0���{�S�͕�%��+�`l�_���<ȆF͝��i���?c~?�pgaz׵4�(�ek����p(�jআ�.3��X��z&��Y1�W��^�|�'G�K��u��T�#
��.��7�8�p�hY�r��Ӟ�l��kY���}�19�o��K�F���OKK9$�I�H�ir�F�Q�Bt9����B/pl3;r���P�ذ�i:�sh��,u4Km�W5�f2���	a�ك��6MF���p,�d4�D����b�N �7$��\I��AK	͡s���%�z��@�6R�Y�'\� �ۡ�� ��Nף�F�,S�ᇺ��H%�t�n&6�������� E�~U��k?���lt0Uw��O�A�b؉p��Z��`���� ���|c����H�[/4�g<%-$��Z��۽��� ��J��0q�\�}2��s&Y�J�����9;M�{.�Dw��8)��$���+�peҭx�UXFȕV3�����f���䡝zc��|���RqP0H����X�~o'F��G|��]���nn��jľ,9!A�������o�}�i1�,dc?�B�="�7��\��H�~�#��d�A	���~�J˝�͉7Y�/��98W0�����c_y����~�{�Me�s)F�Nw|�=+��u͉��>��m��(^IN�=��U��D��F07%�V&Z?{,�ަ�"�{�}¡Ё�b��Oh2��p���j�C���m��RwښIz1�D�f��P�OB����ٜ/���s8����P^����l^ZZ����E)O]#x���`%�ñU&�+�o�uL�i�/�&5�VTS�8�D3#�L,�	Y��b@f����w�]��#I���sO�d!�����C���/��ۦ�V������~�l��gŇge�cā�{��tV<Y�V�S�w��w���LsPN#Efi���TN�]ܹL��v��f�kkKU}*mF�0��U��f�7&Ai���B%���yy#�K_��t�Nu����H��KWV�M�����	�ǭ?�$�6��_�et�A(!9���-"���ʟm;�vK��<1;胵c����!_:��
3R�q\a���d\*_�y�����M��s1�p�&��)�y�@�����`��� � }�V�ʒ��+�~,�A	�����/U9?A���n�_�)�v[���#��HB�^�Ë��_`�"��/�������2�8X��)���֑H��|O�:1�qLD��=��*��L�y����#I�&���X�=0o�J��/;R1s�Nns�fݰtc>z{� g�y�ʌ�3if�ʵi����61z�.����RM�rvN�?=��v0�:�
R�򝟨��T�LJЧ�-�a7�Z���LѨ�D4;�U14�bo�r��"���J�ce4Ɉy�P(~Q�a^�5�i�Ŕ�V<�0��ڸE�� �	�j����3�'�]�_���'��ڜYbh�ᬚ�L�lÏ���"�{)===6F�S�-p+49��>Z� �c�"�\���ߐ̜ۥ^���{��H
[þ��,�}�x��Wf\�n�X1�%�jr\�^ ��G�U
�MwG�Ś�e���Zd���t���Y��G�b�*�=��YqZ5qPkOf�v֮������:z#�{�(i�9at�E7Z%������e",�P����(i����V Q=G vo�
7�+1
�~y��U�Q|M#a�=�l�H�b�ᖞb�ɵN������b�^��Z���eO�wn���T]��#�1��%�@m�C��ʄ ��Ő�U`Im�yۣ�wj���=F��`��� W���\�.��/x8��%nt&ʪ�B�}�R���<*+�o�']I�PB�$���o������lH	����%9��.td"'b���I����ӏ�1�6-�{��9�t��`���wU����@\k�����a�ߘ����}�R��j�_�n5�߻m4=����	�
�w*hg���V��+��^��{\��\�G��lI	:�ؒI w�U�@lXf�3i�[LI�����\5�������a�}���M�/�9��R7V�QV	��$s?μۈ����!��lW���G�3�{�7����×��z�����X~��;��!3V�9�e�p����xL&��ʘ��t2&��ovt���L�Oi�2�c�*� 9����D�9ʈ&F����3U����4?pyT4
`*Ԏ>���]^i��a3�躂�������$�i�eؼ��5� 0�����sS�Y��,G����%Q��mLg�����ͽZߒHQ5�`���ȕ,K�����1F�&	V4`$2��k�}b>�c�+(E?'<�w���6�H�C&u �,P.�SheFDTT����  eS���Q�ۉKk�e�-�}���H(���v�8g��s��̲Y)�L1���~�Z?sR��*�����a (��uۓ�'}R�����OV ˞�]N��;o�/�U�7�V$ �"�I	b�1r�o��1Y�A��:0c��n�5*�hy�4���X�V1�⩵��)�iHd�Q�^�I�ߓ���̦p+���#�ޗ��Gs�#i�x�q�Y�N�r��Y�JP�vCj/��S�Kѵ� �v�8��:�x��t*팊Y�NL��mtT����wT�GN����X�o�J*'��B��R�o��_@t�Z�y�Z-��ksy�6+�G�����4ۗg(=P4W �+�W��/���BG��[viX�r	b�伿h�R?�o�T�'�rB6J�-
�@�$�:}1.��;n�)�L��sC��O���c��~��2�zKׁLw���W��ݶS�<�`���6'׊I$�b���Z����	�b�~�X��)-U^��/�xh��� �۔���"Z��=+|Yȹ���-4L^��*9Mm��6��{���W�� R٦��s�1Ȕ�P���y%F���#���R_�{���Wϼ��87#���G2��S�TDl������X|��E0Mt��}j4�n�����1��6��&�ؤ�<�g���D��矷�c�$�$�Y�Ԥ�+��Bt��)����;����cG0��_�'G")�A��%��"&��_�fv�+X}���ab�:[ؠx�D�&C%/g�dmvfr#�7�i���Ubl�*�Ք��Q�63h��O@i���sr� ?`� -��<d�٪:QvI�L1i����X�]���c�;��o��d	)�i����(O$�>n��({�����ғf�@��+G,��ʧb[o^���g/VD� �W��v�=RAW*Wp�C_��I���TU9�Ҫ���۫���;�}TK�m=�,�BSl��E�"1�"�R�	�iVBƭ�-�%��\�G:@2����q�nx�^�cG�b�\�&l��	��8��r�7;(M?�b�E�v������9�07��V1�J���uoPF�bo$Rj���J�k> �O2ި��0��ĝ����S�H��Y�Lt]���z�pmX `��D���$	�O�(	� ��m~�-jέ9��½�w))��?萇���_��h�{@�j�?�wTS[�.�9�=��5
*D@�[(
"(M��H'���(��
H	(H�^Gz�R�B	=���������q��~�x�=����lϜ{g��L�n�٘�@�/��"�O`m1O�f;Ύ���r�u������b��⽨�g����sV�]tH����_��s�
�8�wY�Q3���,�� 'n�� �'�9,Z�A-��I�
¤F-DےS�����1�}u�s��~���^Ǳ�[�����e�=�F�~y4g��[��۳@ً�>2x��Ϥ��Ҋ���7oR�,��]M�	}��Φ �|�FOR� g��U�ünۣ�����qZsk��h�Ѧ�i��X��-���%��W�1g߸��-�/p�����$����}J��8�G�.������gd�(<A���Z��As�d�X*��*`�1���[�.ݞ �B��#%nv�gά�uH�A�+3��P�k�����O'��&_���A��Km��k#�,0K@wR&�[@6�T�M5�`3�UϽ��D�/���J{HB�4�����Q��n
X K�t`^�k��5�@�t��z0&WU� ��*~�z��η��-{�H��vi%�T����A� Kp�t��8`I�:�f,L��%�3��#~z����aР�����7Dɞ��1��5�>��F�L��=�
h�4~{�·�۝�\e��]^$2��\� o��4	�k�Q �""Co\�2_F3���p97�z���*����C����/��*s��6�B� 1��lړm��5�l�0��(�>�Zl�'�韼��4��L����?���7���Z�1hQ��>����V�0(>�GK0�09������XuE)s� Pf�*�]Qq��d��B3�/:b555s@��1ϳn��8�r��3kޖ�b�20;��9N;��zވ����ϓ�+,%V����Ҋz�,�>��L���B u�dd�D�b��V���`���":�\u���M�� ���|e��b�/�]��$,�6j32tӠ����w�whvM7 ��Қ��R�K�� ���~���~��F
Itն������U���X���s�8v&b���A�H�#Yz���{Z�}�Wu�ں��U�����ҧ����)T�@2(w(,=�7��������n�	�����n� ���#p����Z�L򇒌�n�����f��E��@!&y����DZ�~�/�[ �$� �#ޒ\�;��f+'�35�K�K���`�gN�^�7��n�|B�UM o�ǩ�{E֮��a�c8�����\�`���ӹ��G�֓�������Ѝ�������7�
�V�Bu��7*4���p�hOТɫ �Y6��R����
�'�����I^dg��(C��n��~; �q��H04$D����m��
�22������i����p	��nRgg�+���휢���jv�j�k���z�Y���+����v��[�|�C!�
���Pɚ&S�i���nR׎�����Vf�2���9hw�I�m�#�=���Ô3㪐h]
�4����t. ���`�Qf$���#�`��H���Q�[r�T
9��f1�����/˰�V�r5��>��F/j�6�b1��KQ��E�'��,��95yݺ
:��n�&4�E�8��)u@W^>&�V�H�8�/��K��H�O��+ܕ@���)�[ W��k0n�kǗ�Sv~SWW�i	��uie��{=H�XX���:�_�Q�4��mCG��K�3����L24PK�Ȑ��F���kY�"Bc% ?h��.?��$� !''x*�E�x�q��e!p��&X��7���(�1���R�H��h��eZb��&�u�k���������7��US�K^ML���p5�\ݒ�U�>����S9��A�����3���a�~cZR�Ǐ *w��r����[k�m7F�pC���@����^t�W�hT?{a0�Ǧ�K�KTO[u�qp��m"�: |}@R��Ww&��.&�Fy�P2�)h�͍�"\,������#���PE��
���9��[�<�[�3�x8���3�$����j�Z�-|��w�a�k&˷��jU��hU���{h�<��	-�����$E�!�E���9������n�W���cj�"���$�o���`�c���+�'�*�,q�n���ļ�b��ǧ;d��[�)�+��Y��$G��e�r�����}T� Ց�%�ٱ�.�Pӎ�ã<�f�Vn'�Ww���W�f6]��R�4G�[6~҇�s��vôS�p�
���k�O�V�*~�I�����d�����&�#�.	�6ם*�j� ����Ama�H�eR:�R׋����<��F��
�:�?O����P�AË�T���+5c���-J`��+BI�dS�����Z��<^\8Y��٣��TMM��Tm�	�	;�d��Ŝ£��f�b���@�KPQ����$#u�\mӓ�S�<5#*T�U3��S����%	~>R�)�v����"�����e�x�
i����X��H��v�:i~�@��95j���?�f'����V��S�?̩�7�U���RA��&��El��P�{Y?َ�/?��ѭ�v��j?αRe"�2Q�f?e��(��~�A�U*��l���]��Z�VX������� �����RO�z|h���l����O����Y��N�IkG}ۓ��d�t@B�4g��tm*\�u=��O=������*�����z|CP�e����A�R����T�� ����.�kƹV�hΰ�l�,oY������Й9"��W=*@�z���9X�s*���X�)�-df�����'�/8��T]T��|��|�C�!BǏ���h�����<Ԡ>��u�\l���yúQfX�T�VT�\_� �T!C�8�c�n���>":���S1ڭA��g�����h�.#�1�H�n`�1,�g}��E{��DL������9q� ��
�s0�Q�����tY�\`T�a������OoS�Z�+zJr6xxG']���t��g�l{����UH�+L�Z������I�*.�j�V~���
��R{:��~~���#~�0�,/U
�w��-1��Q����^F���⦵�c�Z��û���=�{�6�� I/&M�;r�1���
�9�FU�&a�<;rgbD�`�1
I��}	d5è���I	��$���}� �����[�f"�|���O݈�n>��DvP��((#�1)��G�����.:�'���-X��,�h�b?�$>����:B���h����8���VE�ߡ2�����Px�45�W#�<��¢�e�6�p�PO&�8� ���;�^`��l{�jFur�P+!@����c�d�=�P����Z�3,}��h�:ի�in���Ɲъ�	��?9�JL���wjO��iL1����O8?��vrN:�9T>4�A�v`�{�^�
��%G�^�ގdo}�\��~c$�]�:���k�j:��tY?��-�zδE���i���s�j��UN�$R�U�A�h�^�0��K���[yB�.K�g0R�lfZb����}�۫7Y����+������L^�d�U�)�E>�\�ں�1r�vB�*��HeJR9�
��/� ���P�.�J[�Ti��j����0	����UV>��m?P�|�����5e���������j�(	+;B��� �S�=i�::_
��H%Q�5,6a�	�Q���ѝ���%ahȥ{;ԩ��An�c�����E	����Y�s�Y�%�Ws%�yb��ˏP�㫏W�OX��/ϗZ�焮�-��.52�ϻ�i�'��w{��-���qH]=�k���Po�G�k�l��'�Sb��\����%�& I��"���,��^�nJSY���'��c��DdA�(�,"ɐ��"��^��C7h��zW45}֍9M��Л����IG���'l��d�u�����4��]C�R�Ϣ����� ���A��$���t"�-S;����,g�SJ)�::}�4���S���m�����B6W�4��K�ȷVb���]�T��9� z1!iE�Mܼ�'��1hj�3I��j��?7�.�F���U*%>�X2 |d+	�g^��]O��O��n���s�ǓHǝی��Ʈ�R�uh�g�I	��3.?I���B�V?'���'����&&s��+d;��kx�9��w����e.�='߂�hC���+����ь�M|���)d
h�2�����/u6_詹4xI-�	k�m�s�]�_���֙T��]��g;�xs ��ޣ�����)��$ �̈XC�3V���.K}Olt{'c����\Nu}�%+�n0#f�?��T϶�̮&�6�s����N�n��,c'�/?���j�D�Y�	�ʯS�����Sོ��"W;��C]a��r)���3T�v��Lk#ߓaO�.�4��tk�u5���(Kܲ]��Qû�e,��Q�q	��N���v��nn����d9�D��\X"�v��Gt�~����X+0�>��mѴ}���Qƃ�.�]��8��'����ﱖy~��.�԰m��ڇb��P��W�9Ƭw�^[5u����SexhZ���Y�Rpj���W��Y|�%�\��(���i���.�����O;�c�s4'��߭ �W3����E(k��a#A�	�D��c޻�K�|A��Z���l�U5:�м�����F���]�f��sgk]m�Cx�H�A�M�������\�b�Y7��D/��k�����~%���z�|M���&��ߩ�Pɪ�����mC49VH�2�$P�HX� ?��=cɯ�q;��koT�<�$u���*�8����J=�؍��,p����)M4�5�~��9�h��C�"9;.,�J�:�[n,	Ȫ�%F"DO�?QcrGN������n(�'�{͓h?}%⁪[F2��y�����$a��sI$~�V[�����������[I�y��E��/M& ШR @hUBB���V�U��_�,ñ��Y}[|`#u��lI!�xϤꣾD����ѵ�1N��B߁�`7�*0b�?)��Q�?���V*Ur��o;������&��6�nx�W������~%���q�r�g����}`$�L}��^|������s��E��}�T5؞��䒗��i٣1bAەx}�E�;����c�B��I!��jHMBI	�q�$�p�݉=>�.G��O
|���9�0���wB�� |��IVRn��1q��O���(��GzSS�ߑ��\Y	'��1e��G��T�Y<3�,�E±g�����S�U�.�����VQ��?�>3=����2�O�I�\��27z/�����퇰��	�I����@tl�}�f�<Y(�$��H���C}���М'bߋ�w���p�l��H|=i!��B�O��JlFT��
���!}a��w^v,�
�����adݷJa���uy��_��yw��3��H���׮�Ɨ�,tܥ���������8��ɲ?]�SD�b��O����'����_���O�	���>���K21雔��[�G L})�_�h�C�K7-#FQ�Bydl����ձI��p���X9r�^A!i�>�&l�󱦻ڇ���[�Kuaj ������\Q�Ln�˱�uhU]��RՀ~ f���c�CjK-L$�б��L������Mu����r�y��8O�� ���0���ϭEWpy�Q�V�p�bg�o��/B��,�<��U���z���L>���P%��/<�`a(���ᾅ��L�p�*Oĸ� �ơkR����O���&Y�W���䩀P��ꌹvP�q]�BR���AgJ7����#�4�'����-	;�0ə��)z��9��f���	9��Y3�k�KmZ���jRީZ��.7���gXQ�a����u1R}}b�"�KY�U)>�_�X�u�b�����KI���d��M��uRO�Їf[khXu� ����">�%6�Ay�$���p��`�t4^������+���]kd�n�x�%6���&�?�����UT R<l�jEz��^���x߷��by�j���O$��|���ގ�	���26e��9���rΑA�_RGC�4��۽/h�U�~��E4N��$�À~�/`\���� �W�ǽ��TE~yPƯ�2��]@������W���
�����(��W]���(�����rH�����ĐT��f�����R�=|.Y��e�,�4��O���8�8)t�Ƈ����+Z[4����ꨁ?>�D$>� Ѡ^��Rkvw�q�i;_
������W^��ii	g���O,V�=��R���Nrs?y355�'��א�]^���%��%4i7W��KUX�g�dgn2ִ��x93W�
K��(��LDڟ�<�V��2�Q�
�A4j�-a�����ȗ*F]�0匈�AnJ}Ή�֔h�[���b�9io rF$�U���yRO����Zݛ	����p���mHn�,�~ms_Q�?���5��ncoxwC����4�Js^�>S���E�l��#�d1L���Uk.U䬭�Ʋ�V�Q������D�����ƿ s�	Y�hzY����
�C��;�I�0Ǔ�g��
�ދ�������_lJoj����+��5{zd���}���w�P�u��/���	�X6r��2���wW&��"z��CS��matt�� _zx<%R"L۴�nҟ/��`�K����~]��y�V�H�v��䮏�q���@����=>vQ1�J�b��"$�6���#9�N�*���9)�IP�1O���	0�wrs��/k�cs��;�]��,V�;;Re�Ml| }(o�oh�2� C��k1�c�`���K��wk5�[��^�4>j�][6��8��t:G�io�f�'�C�Ѽm��t�������3�c͡�𕀋����6ѱ:��W9n`k�p��7�HA�6*ʾw���J��4^�[@re1�������)/�U�~6��s�d�^C.X?�S� 'Yu6�{��=���^ޕ ��u�Nz��b�Pᇔ����^�{��9�����Ǿ���������kJX_$�P�����0�^[�f�pQP9�3*ok���0��FZ�N[����]�C��z����9A:�*��t��>�B!ij���x����<�N��ǎ��l>o�1��\t�����6
��?�����
?Œ:�o���[W^����װ��+'��F�%N^�Zu��k���:����P�6�P��=���K9���
^gx�[V\ҟW��^x�Ԛ�%j�;'���C���q��.����1K�*��o�'8����Ú�>�5)>��$�;��ܧ;3<+����V�2�سp.6�I���w��r;*��DL�(����]��2yz�@:�7ɍ"!���u��U7'�t]fbr�=K���!r[䑳˃��w�>�fhA���j+S�Ǒ�
Φ'[����<�Q�(�<Zc/A� ��8=��Jo�y��J�od�W��%z]ɽ8��3*�w�g͝�F;�2�d����-���t̧]�	:4�QΡ���;��R�&�
e�`��4g(�W�{�&�n�(���F+$&[�m�S�|YA*M�=f���U�D{$wN�*Q��O�Jw�+��o�N��6t	��s�N*M]�o��㩶���#���q��▬z�א�ɻ���Ճɘ>Ҳju�.a�v��me,�=��CD�\���kd�8F,�"�LQ���B4}��6�$���qV.yw��p$���T*�S���䗍mA\�{�`��gP�v��P�L��*q1cl�P����yF��-ʊZ+�sn�+����(5���<Q7��_�H+��C�2*>k�R�Vn�%�r�5U�L��W��ԦV=I_��y��|B*���l���"��Ҡ�B���
��J�>狹i���O��TGcG�v�a�on%j����z1fk���@+���Ɖe�@����������>�&����D�^k��x�3�SIPH�n���NU%��BjОd�p��\`�2�`UP.�u���jP{�]S�N!ӂ�\".N!��Y n��V����=���D$Y�>B�}�>�J3��'��/T�]�KP� M�-0��J�$��<?�K����j!��E���ڞ��^ǭ޻������A�5q����i}���^ͬ�F�|c�f�ω'��Z��w"�Y���:3��h�4m�H.)�R39Y��u�T*Te��ګ�P���T5����<�X �̃Z��$JИ�E#�㳫�����	/�x��-W
�KCJ������{�e�a�����n���y�d���<p���z����f�� �:́0������ �}�D��`���F�PԮ��L>��0D8a�\�y<g��e�h�f��?��T�%|�8�2���5�y�_�VtiB�v�r?6ʀÔ�ѿ��d\��jy���ڟ���ȭ�P6�F+�١>��.�ݥ��;V��%��������
��AC[��I�@[����¶Y�ĳ���t���:�����&]��H�T$��9+(�|muD��Df]�V�]�K����P��>d��0�[֗=�|��ZXi�P:�܊0@8�CM5�=�휎<n�A�x"�:=PT����1��ܪ��	/DfI!
UY;�K��yy��5��W�m��1�3ߑ9N���?�(">��LɫUiA���Q]p*�(T׫�S+ז'������(?���w��K� U�h~�e�.N�6�C�9��K�P���T���p�V��k���vC�|�xC-���;��׳th��K���$^�y8-U�YW��L+o�l;��.�ڪ��J ���o4N%�����7@,����q��~��H��G�s���8Q{����ar��ҭ�ϓ
{Ctdܯ�D&{
���#��/k]p����	;�r�7�@' L_T�Os*#	��K����:���4���.��=�Ჲ���J��k����Wx�e3_8���W�;Aז���m7��@�/�%} ��qA
"��	d��_��d ��m�kc��/�yyｯݬ���f{�#4��´����|_��b�Ԅ���썄6q�&��O�T_*<�{:��I�]��]�yk�
o���Q��8�=t璠��S�ow��w��w�n��~\���!��O]�#*��hq-���8�D�C�G�q|�Og6����v�����@�{�;R�x�lŃ�/L�v"d��S�.<�y���g6f�^1���;�E~A�~�%�s!�#U6^��'�˲����U:)M�u��La�fY���k,vU���:n�5�U�����H!����M6�{A�.j���ƫh�g~F��&�k�	؁����)���˽/���b������o�Y�̚����˫hm��������.9دeIn.�F��oьY�r�Q���T���K�3�2�x�-�oJ�O��)�)h(#MCK�+6j�y��O��h�0�뭱T�w~�%�Ծl_�j��8���'���a��U40�!��ܢ��5�����j��EQn^m��Ŏ�bi��`K��CCǥ[��l���)9oCt��L�L�!�v�4kxa�4ܻ����X1�(�YU<����O�
�^�s�C(JkGjX8��d� �[�)�5jiU����ߓ;�_�7�۰1	��(M�76�4mё_$u\Χ�Q�#�&��"�#��_�LY�_	x�������\+�OϿ,����G=�l�բ���@{��+��c�O t�b���涮S� [��K�L�e��|f��{b�q��$�eڀ,���p��n`���`�
�]�
`t�fփfE��!ǋ���7��ц���:t$��~�;�F��-CMSծ��X������ǊuT�_�c^��I�FXu��b}!ڽI����Yk�VFUD�Fl@��Mٰ���k����)�S��6�����>��ᯜe��i�b*�CV�/]��+Jpu�%م.�ڦ��K�Ӊa�7�M1 �L��g &
0��9�-+��S+��Q�&J��㗍����ߧ%�~m��*@�/D�a�z���"�y\�X2�Ok�fQ��7�jB4�[�s�ۚ2��k�r,��t�usJ>�34b^VuLu-�*y�c��W<tyʪ0d8�`�٫��Ĝ�2�;��{z!n��P���c��Ȩ�o}�]{䊚�h $s|`M�R��i+M�����3}���o�%���=�v�M�iŕ\�SV�>?ZL�oY`D-����k9n뙈zG�k�V4���K>ܫ:`�]����5_��=hC��s�Z�Ɣ�y��ŔX�e�Fs�	pV��0�w=�ۥ�@��Y�SE��a�I�&�i!ǜ����n]KXy>\s�ch2�Ϯ�ޡk�1WL.��5�λ����<@�uE�0�Xpۉ����Fv(,P-�@��".\�����\��ܼ��%�<�X1�W*>�C���f�'�n�߽����<P�{ ��[]&
ľ4���A�[y�XP�Lz��XJ�����fu��2�M(ׅ5�A�8J=��n��{-55����[[�����z�J��Jj5�D��+���P�dQ������h�5����"�a-	6+�"�UHTm���Y�y��u�FS����v��<�b9��=v�ѡ=љv&b�q^�I&MZ�0_ւи���XT��e{��5��aA��>� )͸����V��v��go�jD,�� pH1Z�L3�Y׼l�<@Jս.��`z�*�hJ�I�������|��E�I����`�$���w��ڡ��\<��6���}�غ���sA�'$���!=���2o�|	���95��һ!ȕёb�}��Ux!�f�e#J�}`
�O��+��"�z�N���N�θ^cb�)�|�E����Um٨�[B�"���-��))_����f_�3�漄��w�n�c�,�3�vN�x�(�-Ξ�9�"0��e����F���;7��?F�L1� �6����X�YhO K�Z3!�..LK9���g��A���[Q���|��\�#��,w�H����ۿ��ލ����m�1�}y�mÛ$&��q�q�:��8	Hҹ�j���F#T��⥜r���ue_i���8v+�vt��S��8=�U}#Pu�u0^Г��_-�=��*밼�����N�f���Р].\Oy.h ��s�P�h��W�����Eg7O!�}�>
sk��pZ��#ﵬvg�o�����htg�[�G[�|M8j�9��gby��A��������Қ�Fc8t��3/��U�(��/�X�U�5+�R�ǃ6�>�����N��ɫ�斖� �&ే&��4��@�[4���X�-r��+������Bl4c����	�X(�r|kmߴ��pZ�ޣ�zg:h7��\gem���&GGϜ��v��?9HH�n1]�dV�*�o� � @@���+�Wt9�^L[U�KB3�u�Gvyh��-4Ꮚd�T������Լ;[W�fX�(�ƣ���F�k�z5B�TFUFO"j��#�e���-��`����Y�o|]ׇ@��{����ަ�Ym��
cNIM� p�q{�ln����v�85el�RP��$ �<���u�!d�$���HO��44��o���U��+^����Z֟��;;��ywi&[��m�Kx��G��8��ӗ���R�X�9Yd8�����g竑OX%�D�Fɉ�+�.�T%pY�i�;�4�CT�U4�$|������v琔���J'���ͭ�7?�fЭ#U�x/��-Z�X�Xi$�����v��֭�Ĳ�'�"2J2,Hs��hT��|҅FJNMM�:a}��Q���� �[\\�1Z^�d���ǘ`1�! �o����'���y�I�k��j�f(�Ccs����ZG�J{�YE"i�����%B�9Y��0O�]��J�>mh���y�����`O��4��Y#��xs癱���v�C���9Rr��v:s�Wʶz�z8�N�DI��y���snD��+x!kr��&�Jkh>1���tΜ��7ă��E����өa$>���m8��f!n�����t�Rn;��@���iGb�9K�ݡ�Ϳ�%��l5l�mN
�+/^�F��rZ������4�#��}E'� ��\��&S'��n�y��lN��Z=?�����cY��X��� �IAN=	EW)�G %�BkP����P0�ۤ�u������'@�+�v�lg��*c��F{h�p�{��u/_r�a<ދ)'�X@�I�����U�����]�n�2򜎔�+{W({�N,�Dj����O���B�����H�qJ�4耓�:<@S���f����/^\���Hx �e��ܱ�'-��Íh��H�M����[Z�F�2�۾`�]f.8��m&�ݭO�i�̖>���ѓ��ޝ5�͚ͅ��ꐎ�]��A�ɓ��-�8�=;;�?������*(�/9`@�<]�Y>bٻ����=Z��� 	S�TU���!�:Kĩ�����9`�ڻ���@�oO�VK��v� ٹT�r��g���0��|�j�~v� ��a;��\���.y�,���6��?�`��:__	u�5c�D�G�}���Yt��T�$VC�r�'�F�l螬�[�nS�B)� :�!#%�+��e����� 1�.~��=-�6)z�Mk� 'X�Te=;@�a����	���˫k�x􆕫�{�n�~9����G}��<�6$,�f�	WZ[%��׹��\�^c�z�|�)��S�����x�Hm�����[$]z���Bl��p�R9��x_�sV�Ӥ��i|�]�щ�OZm�[����U�Zz�Ǐ�)�������n�*j�� ����m�R�����66�ݼ���S���Y�s1׳o�QF�s݇6����y{+����)D���s�/+P� �N������K��:^O�A}P���ꀏ�ޯ����޼�]���F��etg����GG�u_u�Qd^YY�zIC���g��� g����.l]�Fo����#����hWӸ��ǝ�;�$��?�S�\O�yVn8Ja2>PefͰ�\e)9�(˸��8�D���j�azz�
�E�-4�Jtn��Q��]��G�"g��$�?�@�s̺���?����/�xu���:8��S���|(ݥ"_�m�qR���	͸���
M��:,�v��3�QA�|���P�4�\4A�h�{�w�;�;j�]�47��.��X�e5�40NْS��U*����΄꥗q//a�XB�lx�X>�O%���|g�@��Y�\��=�{"fD��G�΀bM+�%���W�dS�ʕ�8z-��9Փm
��.mkm�~<��0�1]z�Fd��_��~s�*�#���B'����~��\::���I(W�+X@R
�jWjOAA_�RE�'5�w�*q����Țz���]�%����1M����7��[��s�[>����k�{:2ǄsH;J���"JmO�(W�'O����TSR�HsDڕ6'Q�Hך�Y�5�l.j��$����<:򮾈Nm_������O��T����0�0B:�$��[�E0���r�$�mz�pIIiR&����M���iڙ�~��W?����/ƆC���S����H��%-�)%+�
��K��U�is��ϊZ�X��q۹��&ݬCCC��w��ĳ��?wa��W�{��Z'�1����y��THGW#]��vM$�����6�Ji����
e���T��a(X���E�(�n:0��{P�����+"��g�6���@W�IU8ûg�1ѷ9:e�cf΢+�K�'�6�%"]��띢Lq������Z�H�EHx�؂�u��՛$;}թ���\A�S[>Y�[X��6����' K�t����W����Pz�P�.��T@��������+�,�R����ޑ�\�=׉=3Y�M�w%V�~�gs��Sj��O�Н��W�������X
z}�DA�V��"Q��g9�� �OǦ��s�ͣ��#>�֒���í�'b����{�}/����E�`bo>:|B���ρ�/�k�կ-.oV���SQ�ÿK�K���P�n)�It�P���ĺo<}�)IW�V;$h5m�����z)3��>�۩���C��8��s+XI�5cB�W�*U��/l������ze����k[��Eih�;n�vj���ߕ;Gm�$���-���u>���������s�~��y����p����� �8T"��!���7��?[���}��/�`��g;�9��-���Ō�|��k[;}C���O6�,\��iYJc���x-��j��������龧��U���
u��z.�8���'��p����%˜��`�{��K��-Z�y��ȇ�UznMY^G�&�yl���E�R��X�4���w�·��Α�`�A��8��fjE
t�.�}n��xFz4�������L�NE+��$�W��IC������\�j4>	�e��y�ݬԽ|�`-��1�s�d<������v1A��k��~����xJc�uYɃ�Ur"���%.8��@���90�g�D6]�*"8*Qhl#�����Xln���m�Xf�֩n�k��&���{N���ͫ3+��k&f��>B�&&E+�Sʓ�$�0�$&��(���ǯ����L
SfR�*���H��ERP3+���K�0ԇ^C�� �1'��K�#�MMM�3s���D�&=�i����?�^ЗyB���	�-*2��^]u��}���_��6c)�x���
_oŊ�T����&��X�����Sv�;|�?��W?��ϙ���_���_\��W׽�	IY�MbFb�����{�hZ��Ueܶe=��:G�C�z�d	[�Vcs�,Y;��l9?$
*�?��o�ϗ�����S�[�u�`+׹�\P�ӑ�N���b6�er_a;��#�ݺ�r��5����~��G�D��UV��6�~}��b�
n^e_%멃��4�^��z����Q���E�9� ˮ׆�Q�Ha�Q�K���:g�d���du�/e�׃\�/���[�M�C�V����;����ʾ�eԚmj��%�?Q)J��h�#��O����EM/�(%�J<��[e�ᢰ�֞�׾�*Ŕ�����d��-��?�P�f�i�6j���?�L��ea�fev{}�=������n�3R���y�[���n��kf{O���}3��;3">*D=ݶha<���_��>��9�
�l+((HZ�g�Z��j��>�m�%h�p�6Q��c}y�l׺�5AF�o,�B���#_�yv~�~H���?����vw�:F}�J�@��I��9�^���〇���$����r�٥�s�Qc�%��I����!;'~W0��UDe���ͽĆ��ӓ�QV��
�d#<�'�y3MJ�^�R���t��������}9J94�~�t��#��.��C$�3������g��nf��R�R�G��u�r��9f�F(Ok~.?�!�[oůlp~�������x|C�����Y��.�����=�uO�	������P������'�&�⻬m̈�sQJ�t���ݹ�I;}v?���?��?"�#���H�)zg���ݾpH��jS�1K ��V�P��=Hw�l6�O]1J��He��Z=2���tj���{κ�ǟ��7�v+ܔ-�BW[?��+'I���X��'�׼��>��9f��:�m�Aw|�x2�d.�`V��ĥA�យ�(�@_�%���.��,"�'�o�s�I�;0�[���1�y>�6oQ�U%���.���[�C�t�C�=�[dm��E)��-��#�*{�֖|(�L救�xUS����$�_�P8���[�;���iѩ˧'�Ӷ*ػPiB���'�-�|;�C���-�2��t�`prk��1��@�I�>�C�a~����k}�)om����v����Ob�P��דs�`\MIXw9w��6���#�K����&==�[s@w�,�U�9n0$�V\Μs�ۓ�{�b@1�[��?R�c����*u�OJ꘿��6+�El��۬�=@*W���҈����O����DY��y�Ċ��ʷ�����x�Ͱ{s����F*b�n]�����PtVn�+�9�����Ğ��S��rW���}~E�_�$+Vl{X�\w㪼�����xM��0"Xtu�b'�����z�uM��z��#V�>B��&�:)���ZZ��/<����D,�Dqf�ZJƅ���)��6C*�x�gVz�����Yԛ[������}�oH���=�A�G[/��8u�/�ۓ��ƶ�+������ ��]�|g�*y/�_K'`:�WfV����׉�a��P㇎����e�o����Q�S�R��(�

{����t��-iZny<R|�����Eov&�I�������.M<��6�n"
(i��?���9�����"G�}�[=e�8�Bt1ia�ma8�ͅ��\�F�_�v�z���ˇ�_:n#�O��S��s���Bh�[R��?m��:��o�?NH9!��Meke�ez�2�+6ce&��bg�3⳽��+�Ҍ��R�k�$/���~97��J�����߸�Е�s��L�������MGRz���~���vP�v����������)2A$�ӑ�n�ª����N5����r�����o{׸2�AŻ�I���tmy�O{�<�m-nxm*�#�,%�VUs�u1�_����>��U�V,:��=��ȱ��q,���_2<�"�V��#���#m.d3�:��Y^馻,tt�S�itt��=JV)�r�u��(=5�r>���C#L-����&߭�?�m��KܹKmh'�6,�sN�H����ҝ�m����{\T�Ua���������Gz)��u�D�
�?zq��Um#���N�kV>�g�Pm{%������%ir���b���f���C�|��J���׹�+U�m�v�6�Y�K���N�n%R�+�K��JS���Q����R�Dr,8�'ń�0��e��D�bj�*+	�&��2�������&x/�jdk����ֻU1��7ݼf6�[!�m���z]����C�����_#?��F���Iz�P�ܩ�j��C8vc���-o�EX�EU2}\6cd#"�w�%|�N�ן�������w�W��bB���޽?�;� �N�h��UYZ��������EM� ���թ�����_���AOؔQ���gO�~�wArT���MV,ݫ�W���,��(����<v�O�ɑ/K�w��)����I��E�t'��d4�"u��Q�1(�[hq��/6�ƴ��|���cbC�犍��8{_M�eդnz�L�A�a��� oL�K�.���Zn!��d3�_�(�0������_p�i0��;iӚ�!R�l�6j�༉�uH����ߗ�.���e9���u�%Ň[rž|S���%��~1Օ��{s���kf��sk��P�0aD���2_���/O�}�cYW7�z���J�(���e��K�ߑW���c7>n8��>��;}�|�G�]���;��.�[��O�������?��
�E'I�$9v)G�.��f�k�<u� �[Ju���q������Ys�VT�[H�Sf�to��i�P��/�9'Y��K��Ysi2�r���ٔ�]=rcX�.�9�)�\�L3BL��?��;���}���bAQ�bDE�"$4E�w�
� %��F���HPZ��!�"EP�z�PB�3W ��;��s�8����1₵�|��>�\s��|{f1��xx�3�|��x���3|O�iG�B�8�m���r�'�H�PG�ʱ۞�.I��Q��W�?�[+�&�Rb�`��+%�rK�x��}�_��.)ﯖ�A�9tj�̂肏�F㵂��y����1�4���O�,�J/.b�H�btuS\�\r�aolұ�q�艜�������`0U�T]R����R��N`�!���	�g�	i��jfƹHV_�6:�]~��z�3�2�g��GI nqR�#�Qg�2��C�2c�b���u
�eA
'��U4���eϸ-'|����E��+������?��/�k�?�D*c��[����ѥ���c�u=�Y���R���C�t� ��4���7$Q��J]Ӏ�6��)&a?]�d��`e�%/��.g�5fae�Dc,G+��~!A�2	-I�����r��������hJCʺYp����C��o�S��U�I�A�J C�E�^��/¨p�˅�.��u`��**P ?"z�/-2s!�y_���qE���ɶ��aݜoB��:bhQO֍�ṷ�A)�S��"����,�E4��;5�;Yr{�������dN$r��<� �%���K�i���N6d��w�}��x;�޹v�J)�Oo��q���h���~e4�P3��� 1�;PhL���F�j7�$Иk�loT�h(&�Ԥ���}O�g�ꨪ+��} ؑ���I��Q&��Oe犥���bG�mV���w4R���]꩞H��p,~;���q9����O]3^����R6���i@��<r�y��,�RW�
����:������G�{�vkn@�}8���*d�G��%t�[M4���0���xO{��<�IYf���#RE��u)�O�2��Q��o4�尿�%6�#�֭���>HJ�����
I/m����s�ט�s�1ӑ�|"D�U�˺
��(n�TF�7]��`���N�z�7i(���Sq�ֵs���X��҃���׿���{�K��K//,g�:j�1y` h��/��r4K�r�PM���m4~Fc�GISQF�㸨kB:�}�;�/@)ʛ��&fd��0����e�
�**ǷL��{+���x��8�h,,sA�=Sc;i�����#�&����J�W����#��U��0���n�y��V���N��w`x��6&��p#�i��z��<����*oi�o���_�w�_4A=������>"�^{��/vG���/���b_!����M`����+a�]��_Oz_��y��"�]�Sxy��G�������'"�Ul~3:!��+0rCc��R�N�7�r�/�T�r�&���T�괛�~��0����C�J�h�oZ�l��w�,��/���2χ�p�ع]��E��^��jcS��jR[ӄ�9�lK 6��.GT�l����v�1�N���R�g��չ̸��	 �_t�U�����,�7��Td�{�zg�#y�0���S��7�_���o�8�
���� �h�W����<弴�Y�R4kP�h����@f	D��=IIzq�ɋ#�_�P����6��2��
���W]����_��7�t�C�7�u��+�h����;�N�dN��?����@���F䩈Aޱ/���������|�f�ς��l��3B��~�ȋ!(�v�<[�D�n���AvW�/{��V�W����@C�<��y:C�3Q�2
�Q�"�So���=Gt�ܗ��2B���Z.��� T}����B����&�<��V��";��?c�4� �bW�]Ruv��Ի)��������ޓZ���IR�h"��g��^��?P���Q�ʗ�O����o�� 1���"R�_d����q�S�i�uɢ�{������N~�}�"�Z�X��W��u�Cc����{��-C��9�2ۍ�OǈK�e��}��\ 
�l�'/*ۊ�ك��w���&(G��[H�u�t���Ŧy�{�L�by��,���b��x�\�jSE*u�Rn��
��xI1������}"쾖@�U"r����A�=R0D�X��M/�$R���ݳ+ٓ 8�d[��d[j�}����#��T��^`ey�1(&!����9��2�H>Ewz��X�-M�tK����Oɇ����d��LN_p�Zv���v�nn!��ñ���^	��J �@a��Δj/�Z�V��j��8�~.]?���:�V$���)�Y3�l�a@Nk��$�r�z�a |Dws��zv��r�cs�g�
��oQ��J!3���K��+g���Q�]���oZ�[{�� ����{���M�s��|��\'~�݄v��'�Jy(����Uc��e���i����_db��B!�;sW�{�v���x����5�aU��2�}�&������Pz˩��� ����۾*oh�]{p�co��z?
�;��IC=�	��	������ {����Z7
�Fr��뤘'Lh	����fC .c�DQB�Tcm�'����'N[�LD%&���
SĔo{��k��>�9=�0u��JWJ�eI��=��z}@����Hr��Ձ
5��8��c����4�c�/,J5�A	wk�����Gd��9���� 
�Ի/�%�@q����2t��=�󏦅����f�8��Hl�&��n��.OWX���s]UV��^���9�z�z��~�F%����IK�}�d��	�P	es��/��L��d�We)\5�z�v�ґ��´�c�A��� k���<���~�W�����Ꙏ�f4�9�1]�$}��c���p�ƲT��I��|B�k�YM}�༃"r��ɀҁ�a}�""wc�7H�p�KzQV���9z?��(��joi�΍�sW�f�%,�N����j��O�I��O��������)M?D'��y�c'�ͩ�s*\ Ƹ���>�'?�t���2��H�G�$c� ()p~�N��V��`nc�R'�3��D��$��k�P��^���&&�EJ%��CH5�%�V��ӡ�E��c1Ά�٠���2=���%ÅrdJ�����3���)t\��C�Q���8 ���a�,� X~��^�@v=�
�����f���I{�}��D���o�L�\��P�#f}����9-�EG�c>����� 9ʋD�E׹�nD��3�c׻�
P��j�~�X_��sP�*��!��YU&25aL��r�eD"���~�U���鹯S3�p<���P-w� ���~�������(��Oɇ�k��U��:��C�~%�L�0������2�������N]��<�i-�9��;ya��94%]�.2 ���D���P��r�Ʊ�etN�S��q�Zɮ?�Ez6�����9�
����6��b�'2�_��������+kH���|�5!k��hV�xƧ(Ue����S9��MO�Q2wUYbV�T�2�k[�[���R�90�Ѡ0��P�~-�v�&c?�ߐ:U1<�-�8��*��$W2*ZΌ��9�
��.�k�������w��Y��M& #D�¥,��q_�^e���2c�s?\��4�?`��\$x+h��Ty��/��6�I�"��Y�5w��D]�8И���}���l��Z����}+���Uf9v%�����2ФQ��̔�0��t�:TT�,���h)[������=�y��c�� v�����QM{~�h�KLKoG�P����*ui��T��lU����ʎ'z�]�0��0J��B����Ť����ZǤ(DJy���a���)��RoM�o�w��(gP�U�6W�5bC�ث�XȰY�m��</�ܷ�:�O�z�NS���ې�Y�g�B�QPR-lK�Bi��Z'��z�=�r�3V6���V]���\Ա�C�y��!�fI���kH��>j��o�u�#�4az-	���p)�\�ei����V�5��O'����eȞ�Ъ�������.��	��������d=Lο�x��2��i��/�����	*.�������IJ�\�K	�bD��N(��N_֡��U��!+%=�f�k �m炱����B�0hԠ��Y#,{�]��4�0\ )wx�������^�Ѓ�fZrHx�*S�e�kŞ䰃,�Z�P�s1!mǷ��g�Hر��1�����PL�޺LN��R+A�R�a�� ����s��`��g�����z2���"�-�afy�bh��,�o�h�YZ��b.��]��{����x�1��k��0�3;@�n��FOf到� ��v���W�86jy�I-;�3����~����g8��������8k����+��_9��_�=���Y��|�H5��=;�n�SX�����dGt����i5�@8�Ж�ިX���g}�캈��h�R|����E��J/� y=V���aĮܵ���x�=���y:4?�T��O�����kǎ�[x��Ž1���pw_:�q6	�迓���#��]��ݗf��&��IE����^���B�aMK0D�#K���2�1�k0�ٔ�A_U4sb�U��*6��M%BW����Y�4N�.�	���m�_�b+��q_Ķ\pq|�N�Ǿ菮��z�T�.�	������ݴ&�UO��k�=�_�AEu꿪x��%�P�,s���$�p�y�E��V�0�oe�b�oPm	��v��?Έ��V����^e���:�������%��5���8sC\@�L�\�t·\v�1�|j���>ij)�`>W+���`�k�D��-S\%����M��eC�)���c�x��%���Fn���R,'���a��-�`v�#�3}��3Z\�Gk�e1�a�l����gT����>���q��n�x�

	1��{�3�{�]��9{K��	�@��
���M��O�/L���M���ύl�.E�bS�� �H���9jQKDJ�ne�U_NX�}��2����cc�����r�r1b	X^^.~2��>T���=��ʵ�\����L�ݯo�-T�DˊM��ފ�^i��&���\�Da�'A�$K2u���mֶJ��-12&&��1�7���/e`��?�>�S�e�Q�Y�U�V��%8�_z�1�����U�|T���ux7,���������j�F�WB����E�����OK�������?��?��������g�حm����g2+��8���#(�+1-�H��8>B�B�UB��2�hהPB��3����19�E�;����}E�7>yO�R;w/]�'���K��h���>�\}�v����/ND���(�r�4��R��r�N$C���T �m,|��v���R4L���фM�:�>~�����7ω�4�q��n(.�֣[���պz}���Ob��w�-g٤�c�����Xf��q��J�i������=�!�����tg�;�����A��c�l��y`�]e�R/:`\k"YT�|hX�/B̈́4�����jω���Z���m���&�ض�����[Ô��ݯ���z����ve*�'�w�^,����N,�~�{���AW~���� ������OĖܓ;Q��ЉC�.3�/�+�lj��1�ؖ2<����A%�/����Z�~A|e8�D��LWqZ-�y+���Q��/�1����Au�:_9�3�!9{�b�d����婱�@�lG��n�
��7;r;���Z�IԾGl,3�H��?�!���O�C��Y��Í�oO0hL5m��~T혐�|�5�nT��q�[�����YY��l����O��}�6���t@��O�Z���P o�����g����gr��i��ӟ�n�?���D_/ ���D���zg�Z�idzD�/�u&�/�:?��Ոsē�����hr�,q���y�c���αo�ln����fb�����;�����XqJ�L��?��`4�_�@%�_��������m?�%�
*^
lGh��[�T/��}�_-t-|��x��2ڸ(��Mb���r�����OxiA��s��M�:�G	��ߓ�
:���mL�IO�{�I�?H��tR��
�6Z�G�s�	�Lm2#aY`s^��C�6�i�Gy;����U|��γ��Y$K�����6�j�=��Or~�/�����S���%s�hFOX����c���x� U�����?��g��I1�4g,;�K��#��05�՜)�To�"B{Y��Gzs3j�ú�?��[�6�u�]�Y�9����Ũ�a?���me�]]��94�9܅F-�B_��h\_����G東/_'�i�[�x�)�rn�Mͻ�r�X�2�4�q��%�/�f�y�jH�"�Mz�
J���l������lR��_�=6�茺5i&g�LB*uCg��0�&D�hY�S��l}��VA@��D����>�ͥ@���T~s�}��މ�tx���p���q�!�R�٩7Ʉ��J�7���n�Ն��S�~��8��aR������m֬�b�~&E�����rq�g�C���}u�W�j&j�O�;��D������zr��o��H�(�|������il�;�-��}��w�D�i�X��,���W��mwB�ܜ1�9e��[�^�h��蟏$�k&
g��YD��X�"��q���18�z�@,��▓4�E���܉K��uV�T���N;-f��f��oC��IO��[>�+�a�t����U��iA�D�[E[��jh��ƣ�ԋ,/w�寐BZ����GJ�5z[��>�TR�r�i�U�>6�1E��ǳ��(���כd�:�)'a�J�V��s��jN!	��:{!h`k�x�$
��"U�m�ơh.[V��X����ΚM
:f v�����rS��6���w�-ھ�/[�/jJ.1�GJw6L�R�RUWf�T���6�����X��u��<�����T�9����XB�2�Gٙ��؅Q�U��
$� ��7����@ qY�l��/o%�D�P����X~�Dw��h��w}"(�q�\ջ+n��-HǋhLfxv $?��Й���D����1��Fev���.L̀��A�,�!�����=>,b��AO�Z:c��}�M�^��1+�U�ՙ[�RE��g��ތ�~vS��[��T���7J��l��.���fqȷ�2-*�iRC�{�i�1�������8��<��Д+_�v�E'!�A,���e���ȎL`�J�\���5f�¯����/t1�?�R_+��+"�2�7�s`�ki��}u�.��.��K�b>+e|���&}[�h����V@�א�p՜�	����.x��z����i��&_��\�n =��.Q¯�1�OCe6�}6]l�A����ͨ<�d��1�p���bS��u��	;�kS����������������W�1���mX#'�`�r,����Q!Ĉ	{�W��Ȱ��.�)�$ljz�˗��y��S��l���1{(a|╰f��w����ܛ�3�p���~l(�rK��)��N�l�mձ�K������R�h�3�`��a�����U�rub��0�!�O�+%��}�̊.ݠ��B��[�(�F��(Lz/�n��T��2'���Phk��$ ˽����!�n�ܯ5"Ν�fLpXq$º͙�ax��v��ծ�~�|�V�9òc��'?(��
ԭ̱�*�8N���6l)�=9�B�0>=9�3H�V�R?�z�%�K5s$7΃�I�B�fj���V�N=���L,raAӼ�
�x�a#S��
����q�Hi��Չ���߀p�Kq��#?��vm��LX]���=ej��bi�l�N8l�ϕ}�q|8&|[�?H�Ŧ�G�N=#�A�Y,�OK�u�x��ᤸa*���?�"�mH<�m�s$�)��9�ߑE7�����B�Y��S>��?ĝn�-��A|�O��r�>!�dN�L��?�^�<�t�#m�G~(\�+�E�x<�~.�<{Ǳ)��K��O :?T"}D���p�\��y�q�T�o���ʛ�ג����shu�W�'U�s������5K��<h�}[sL¸T���hB�Z(���N�D��Q���T�N
hξs��s���/��;�&��^�}�Z�a���3̨�o��=�L�
�{ç�*���۱Ŗ<�u�����%�MTM�Z=�g�4�!W�P�)S"z��H�{^ϓg���1,ŚI��'ɩeia���nB�v�-_�<��T;* �}�#�M���͒ח�}�?�Iռn& ��>����4P.4��h��@I�![w��9���^�`��_CD�uޖ�~��70� ��!&�2���k��}!�~�I>C��᛫��gyv�D��I�q����m���[y�ՒϮ.f��5ka9�,%��t���x��(0��C�*+",��=����0CW� "Ӫ��ݮ�����Ge�Y���q|��g�A=\v6݋���N��<cm�RۺN�ٳ��)C�pͺAݞ ���[�V���S��N�!�~����e��_�a����>���z`�WW�+
d�C��!���~����%��� f�VG�(�Wˤ$�/
O�2.f���V��W��}�k�Eԏ���UgD:n@��a��~:���6h�ϯk�GuZ╎��t5�T,Tcy��������Q���m����=k��4��9q�*3�_H��q��c;��٦��,m����(�
�|,s���e�
����2��X8�0H��Ɉ�KHƦd ��jvSVU�G~���CZ��eXE���@U�{ٔԫdP��<��~}
��k�V�釟����d�3�|{��{
��?��x��ti�o�l9��3{����̏���R��vp�,�Cy��#�\��{���6�e&ˇN}�ed�춭t��.��u�6�K�N�4 ^�*fTw���U��u�詚��)�*���<�s�����F5Mҵ�܈ j�-;�h��~	�OR۔T�)'������Q�khL����"#7M�u���Hi�ڹ'c��=+:?��z����U��Po����.)��ʵ3�<�<j;=%�Z���+�P8hFup˼<o*1��$�q�*plUPFZf4M���j�,q ��26�b�+�@�a��[~ئ�c�m�U�R_?tt������c��!LB��9h�D��je.�!����%���-����M�����{��t\��V3�j�S#{�'�v�5G�<�> ��u�%=K'N@�o��^�_��&�9�>҅R���x���B�js�04���O��@qҫ��Ɠ���J����7��Ep����	��HY�\�j��Wq�^��_�����|�ٜEZGvu�^�yڻ=���4���Z��[Ъ�w������D�� e᱊�=%N~)���zji,(�~�N�t.4�G��M4����|�\8�$�VR*�f$9LX���:�4�0���Dn���R~���B{_��̰�� 8Pc������:fͣtU��NUULps��(�|��w�`��[|�!%���~��aA�p
���΋nE��[l t�cU��׹�;��ih+�y�@�����N��[~qPϥeY≰��
�8�Yc�$&�؜�9�kj�2�K�O�SP?���T��C��'P;�sD�1G�n�QiIr+�cU.�B.,'���uU����nb�\\Z*r�� �Oi���
h��0[���Pă���WI)����F�4`�n���L��Oƿ}�t#!ͧц��}l!����Ufc����^m_��Q�����@���� D[�N����#A4M�-RO�Y��7`yO��D��(���6�-�F���HbR��|b����
��+��g �,K��:8p}����7?��0��]˩MGa&cu��Ft(�j�䇞������qL�ӝ�t�ya���d��V�`lh����Vg/=�́��$(���= ���2X�k�o�)P6��ޠ�7i�-�+>�ϧ��a��o�.�����Y�i�����R�U�Olŵ�N@�kG���0Az�^(����XE���?��zS~+v*�j()&e�(�A�����nn!�>��j*)0#�s������a7�x� ������̉����[��eC�I�xq�T-SIY�崩c������;fR����sm>۔H_zo��_`u@_D������Ƣyކ6�QfH��޸��TS��|#띺ܹjt[~�o�Y�R
�Nu
a�Tj�� ����K.q�w�&��粼(��p�N��O'� ��Le�'˾ڔ���eϦe[��������#ݓ��Y�t�UieP�t~�'_�B�B�S������	x}z��)�U�8i�Nd(h΀
1������sQ3U/��"ʽ�L^�d�7�K��(����˄���&#�� 7��m�g=ס6��^*����`>��
��V�9�̷���&/ٿ�![��[��w�!:	���t��ƚi5I\4�E�9����d�n���$�'�ʗ:Y�bퟺ1�l��5�y��ħl���˻4�JW!UNZm�mu�?�� �(�JV�Rp8�#'\
��,�6��Hf�SF���x��]Cg�����R��*hIjK�Z�̰N�W�@�I�z̷�H�b�⍟�V	+Q�-�e/��U��g�������;�H'��e^ӱa� �i uK�_�~�B�H�y4��{�y��� ?�q./�u�_[e#�R�#`:�E�|�a+�~^�R�@4���� �D�=:�WPc�Ҕ���ضP�y�TA��n�h�S���a�qu�t˝�*m7��N�\:䷥d���+J�C�Pa�*\I:tM��.9�y��r��ko��	iG�^�7�w�N"�ԏ����}f��j�Y,4Pz�3`��A/��m�
����ގ�� ubL摫OK�q�dq�J�CT�/$玲����Mb�g���
͡�YR��/���/mTd`7�n��d��xP�)Q�W���ؐ�wo�����9ض�\ ���wS�:Xji%ᤲ�X��-C��wÌ�:�e��U(߁����%�?��#�y�iׅB�� G�Β��|�`��T�TGR2�{��j�-���`�h����:��ȧ�.���C������P�˗�׍���}�~��xt|l�Y�9���c�!L�cIs�Ҳ0�;�[��2���4��������gQ�����s��1G���D��>MR��۱9LS��`����f�|���	�Lʓ�UG;��;@�q^�4����w�|��+I�.�Ѧ`'�ZͰ�g���$@,PXn#�-��蠖H��	b�:�[H�}��^���pQ6��������G9�w�*�`{3yh��^+�8)����l�.����/�a)\�]�*�1���'��h�i�A�SM�X� �vt�@�%�k)fa�Fux�kt"1?1�u��pV��Η'���Ql{�Vڷ6^�&�B�[����g����+�F��}w'���	e��*�~ЌY�5������z�Wf1�uy�E��s���?��6���XB:���  �uA+���7�����+G�T��a�J�+69��y���!*�ѽ���I�J�Of�a(�\"�͡�&q��F�p��>}�jf�H���|�18U��DfbOl���1�(A�H�����V69�G�����k9���?�mh3����~�� �R�zM��	� x�k ����@����GuѺO�D2t��m�8k�t��mщT�Ԏ,�p����5ӎ�<�mX�ba��6tT`��J$r�v7M�(��m����"�:�����u�a�2��{�tSt�|"6����EM���9�-s�3��lE�+����P�],��=��@�%��e0Q:�~gށVtr�i_�IKmQ�̪�C���OȌ6"o������X�uF�zeB\N��G�D#�c�V�|�S�C��m�'��P�'���7��u�C�2T]�)�~yX�R��ab�x#A�Y�؄�����Ne���Z�.����8��?М~�m�8�?���:�їc\�r���\V
�إ��	�5�^���m\v÷#4�_	�Eԍ5	�Z`i9�G�Q�I����t�o��d\�i�
k�C�����b��M�iuI7@���8?�*g)�<u�����6�p��G���<=�� 4xg�ywM5��%7��4ԋ�1�(���)tnO%8�d���d�l`<�d�4��!�;"-e^bh�:W�s��۔3�h�e.�L���������!��LN�*u_r�oR#����z�9  �(��r����<���Dv"��)k���~ꑺ6����PE;�Qr����q��L!�ۏ���Ay���H��A_�)��&�l��w����I�M'���PQ��f��\�XN@o[��<�
��.����"JіD����bX��:�`}�n�+����.wծ����"I��m�0��®pZ`�u'�8ծ�i%1�+�[�'�@-C�Z�����e<�T8�1E����X�����]��u�4�P"�!M��k�����{�n�]f�	��ֱn��ׯ�Y��"�*�>���6Ƈ��D >x:�tbLї&����A�8>���gh��vf$�j�����itYQ�ϙC꼶�F?�zkZu�r��Nӳak��k��,����d����v�h�"���{u��bϽ��������Q���!�����Yi�)����~�l(�ӛP�[�"��[lr�Cy/�F�+ؤ��6�sJ���;vN�Ilz�ne����U����[�	�[V��)��#�ޛ�ei}NQ���B���\"m}zNw���`�Ƥˢ��ո����>{w�/�� �,�J��]����C6vLUp�p��A�z��ą����^[T]F���ͣ�S�M7J+��T
+3������p���u�t[	���|agjG�|Lh��{С��xoa]��"�J�Do������;9�<۽]󳶞�Kȡ;;���.��z�ۄm������UO�DR���[_p��\��Z��љ�3c�*S>�XyjtU�É�Z!��|sɃЯ��<�1#����L%�Q���Ȧ�iR<�@n��uwJ���V��t7�dt}�v'�(u���3���;ەߘ���LUn1宧�����26����W��Q��"�s2���x�׈�	qƽ���e\������7������l���;}T���,L�_���ᰲՊv�<���u��u���JHZ���S�Q������."�]�FK}Ɯ���P�C�%��35�V��#�(Ƕ�ve��ں����%j�T��o�������\�C���$Of���=�2Bݠ���PO#)�z8i���D������X��Z�&$c�������V�����6�,옍�0��U
8�57ֳ��?��N�� +�-��	��4��R��l����`�/(�mU��6/"	d~�ݾ%��rw�왱6@ҫ���L-���B�͔�jM�F��ׄ�˼�ݎ�'��]{IR�5�xam�Ys�4���͢j���3H2� S�6���p��[n�J�B���sl{`�6�9r�J�-11��EҚ/\\q�1�u���C?{��pS
�xr��7_-����dn.	Ҙ���U�8/�:�l'��d��U�Fw�er��J���?��يl��P&}b	��YX%i���fz�,�������.������Y3�sU�%�>�j7��Hh5W~'6�)��Kuh
�N&�����{/M������C�2�"����PE#��=i(����b�d��W�Z��/kG���
�9+9�a���H/�����*Z@d�즐�v╽�PDy��/�a��5s���m7(&)�!SAz��wy/_����{g�=�	\X��e5�xA~�Qw�S�����O��p��`�����B#oV�V��R-����(3�읜��EE�{+�z��Ā|��k]WT.��ӧ��k,ct@b~���g�WPA���m��/ވ�����Z�T����mb�h�lx��3�:��*v���6"�s&
�bǆ�C��Y����f��}��F(�v��v���{����,�������|�SKcoίz_o"G>I���5��хNc�Cw��0	�bAm՟_�����$h�[Fr��{�MB�i�oVlͷ#,p��w#�h,���<c���H���x��M�}���]~�z~�e��>�@��;�>&3�k�u��T*f�bt�^�#�xv��b����bE~z<�O�©e��"���Y[oM�F~��˸�j2VY��N�bMx��l�Wmkh�Dm���p���� ��!��{a4僥}� g��Pg��j��)^�b32�a��w�t��M�03q',HLL	H�\[b:�h(��zR\���;}LS1�b�Cp�U��\Ut�bݤ�B��EU��:͖�kQ������5�e
����?`���S����8(�<BV����C���ǝ�z�d�5���&_��	�t|4�łH���f�Ά&^��k���U"~� Շ���X�ʅc��i���Z���i��Z�R�\�f�g�]�>��O�~0hEsg�ě\ߦ��S��Z����A�]fD��h��������o�����d|ǔT1���H�7p���b^����_���$��SS�$;��,���v��ɤ��G/s�=;��t���,�<zVP>=�J��Z~������1{�yܻ�4�VyGւ�|"�J��lqo�� ���.��Ü'�Տ�ֹ����]�h�i�������4{�Dp8�Z�<]b���.{y��1j�����F(��T4O�d�3u���s���%w/��L��ֳ����[u�\x�����m��*���C�pYp4��gB��](�B�?�t��C�y5%6���0��чt���a����db�QgT<F-�쮍58ii[�&����o��H?;ĪE$����TX�73����l��ɴ�W�V쁪�����O�|����:�6j#�V����4�Q��9�{�j%S��Vl܉=�(��j_|�x�VO�P�G�feK�_MGy�q\��3o�.���"����Q[��j+q�W���ZU�S�	�^��M�"ի��{�T�c�3��������	sKn��%�BP����+{.�	��4�ύD�L�<���CΕ`x��^����Jr�};��reIƄwO@��{6�v�R�G���-��>���*6#��u�c�=��c {�̈Ǎ=���}u��Խ�z�����tͭy���t�׌�ߒ{�T����,��kW�����T���C�aIIg�Z��s�$[X�b��tv*+�qB"M<ͯ����V,�OTfK~ݻޟ��z��N�ŊE�CJpe��(�̱�/HL�O������O'�[/.��҆���+h���nqOav�#a��rۍo�zgg�MMz<Ή������e�(w���4���UT$�Z9�nʾ�C�Gk��:*vRC�/��n�?aR=���>s�����1pS������ݕ��<�g������;	�rm��%,���K*	���J��mX*�w�Rǂ^�q�����R޸�{�<EH�H�����7�[s;Kh�tW�?q�O��C��'G�W���Sy�t�k�z>lq�A����Yk����,�]�)�\�1��D���z4�%N�$���m�m�$�A���x<8��m�Ɍ�ʔ	14�i�3���?��pp+w��碌@��X��t��\�{$��Q���wf���obΥJ�=Z�z�)�!�d���ѶB3C9��g�#ḡog��cd_S>��'��w���n��dvv� C�m��%=@���R5X%�ٕ����=9�E�ШV(��=�� ����+g�Sc�b��+��.���-a�x{y��.��ɟ�:��Qm�'r�#5=+�V��l�H�(���@�ѮԨ%��m�b���ߥf��W	䳦W64
eu,��Us�7/rsSc�WGƍ�����,8_4.�p��G�%҆��~��9��6>��,R %`���]N�V�F��HA`��Q�8��~s���ߝk۵�Ru��A��k���q1N����5ImX$hv\��uD��ԑV�_�2a�ۺ�I�Iw�32���L���x3��H6��������2ȣ[c���~ye���`Hp7󺣜q- =Ȓ9>s�zH�t6~&E˹.�%��Ҩ/c�U�E5V^D�a��u���N�K�7�Y������3�w9þ��ߔ�u���C���2w�c���]�fK�J��Dk�oV���n�i��v����g�I�춳��H[����<����2h��>����*_��r!��˜=�}��k���?�Lx>?r1w�A=�*f�]�i��+���?��Z�j-=�[��6[K�s�ۿ�'*$�{��J4���T�Hx�i��写��v;xs�G��3P�9l����+��C!���^G+�y��Q��!�2yZj0�M{��$�==Á� ��߁�T�&���|��kC����'��S����Tڸ��"^zjB��@��i�u u�$En5U���� "Pu2-o=��������g�j��M��*[�6���l`�Qj� �Cc��^��/�昑(�v��S�d2Q�U�wa���ϿjP�i�`��HÇ֍j��Q�G��fY�zZ�R�(-3��8�xX���tQ��B��k�{�U%�iq�7z��Bh��g
���o������k= �u�Qc��S��4�� �c�0AN�5W�� Yz5�g�T5h$���h4bq�d���1Z��%z��i.c�:�uC&���Dzz$�E�`�߾g���4�?�l��w�]�o�@���/fkeU�{�yL��['G�5`ԅBCӞ3�8a��,W��9�$0�W^	|3���E�7���8ػmX�����[��ڰ��'��e@@ ������3�,gf�dV[k�HQq���y��� �[g�A�l�XU����6�:��_�Pb�3��k�g��[���D��p��o�NlPU<ن��](;g̾a�g`<Ei,q��?c�� Y�م�V�@^e
Xy��Z* WZT�4�[�!~����O S({�po2�}��bD0��J��CO��Ae�laV�"�so�JBl��U"�%��b�-+�6%�/��j�\d�ӳ���t��3�����_����D��� �Yx�0˝��]	�R���m��R���᠒-��������w���V��yk��-o���Ox���ڊ��a��QU�E�'��oC(��v����RjB�v�?���#��x'�Wa�\mљ���e ,W1X�Y.彏�Y��I�f��XE��͞�tW��RgU]
*���|o����w��N��j�g�-�H�:���'���=�_W�MX�i��sת�ً1VQ\c).��K���[��rwm��_\�k�[D����$~}�������H}�3+�K't>�O��a=l������.=UyA�	Ya��tSt�R��Y�;W���[4�&ZՠǛ��)�	���cr�@ݻ?ݑ���ͯiX����$���=Y
���^�q�]c�����>7v�����y�Q�J7�E������?S�-�^���B���]�M,m+��F�+A��[�].N����ȯwIow|(�Di��@Ttt��ґ����:�+��=P�L$�H'�!����莧h��A^�۩�yս���/횑S�w�Q�R��bc Nʘ�3���P�j�rϒ"��X��R���?�s�h
Ι�Ӯ���[}�;)����5@���6�m��2�$����r�������z��Ǳ@���.E�Ai�IEB	)I�R�F:d��iF:��r�{�{��������7�f-����>{��y�9 �-�Ij�_����a� Z�f�4͉����[#�7��P;���;��:s,R���X���l V������~O��߷�����x.�l�&��9�����=;���JBݟ�7�V]�MD�Ql�ت�Ab`�̭-�7M�R��E�e�?.��v������`��\%��$iq�&h�|0��a��u�g�ڨ��9��T4���aK��`�����cqNx{U��[�ۚ>����?���&[1zQ�����h��A��I�V����D<b��_ ���e�� �1:�_���Z/&�)�u��2�!��������{��b���,&99��'��쭿{V:Ŭd���G��z�g�P�8������b��	�8Ku����q�Q�fc�ȉVq`�7�Ȫ^�>�4a�IV��l9��ut�B��Q��v(_��q���ܼAn^`'N�S��4��4��-����ku9�Ȳ�����S�p&1��*V�����J�V�Pkh�㟡��n��hۼ*e
��#_��UW��a*����3�0�еd��"�c�q�?"��Ā�6��x�:�3���'�q��A����X�ٕ��y�Zt[�hQX`7�[��nC\S�2��ە���N?��+Z!ۊ;$$@(�w�}�`R�X�Qj�;��=(�=:v��(�Q#FGk�a(�sjx��֢������HL65�I�-j5��N���̠�%J,����ϛ6r���ѡ�%^H�6�Mq�޼���1��6���H{Nɖ@U`��"���NL&|��2{�Y����G=�c�!^�S�F�<��(*�[re🡶���,��Q�����p}u�ͳ��N
�w�~|�ڋn�j���,�j�Np�*�S��o�KY��fS���u�T6�#w��wvܷ�I��ȑ�i(��Z�<�0�'��7l^M����]]�'�z2�O9h���\��0�k#d�R������fqUR�,j����ΆoT>���I�D�ƒAm4f��$�V9)��f�j�=��A�vo�Ǘ���O���5�Z��<�\¤�&z���/F��V��h��9��	�Ye��Q7,h�VreG��  2Z⇇�
q�_�
n����#��gf���'�P���hB@㝂�Ҟ��ő�X��Mݡ*�7v{�l����dY����WQ/����ɓ	V�����"�r����w]�O���;�J���v�L].������կ�2c���X
L�ťƄ���5���u謪��@��|0��B����?�T���7��
8��#����^`}�شN�8�a��'�����B���'#E�/vuJ~���+޼���hމ�IIv������e	U๕����a�ǍU�A�#L�&j���,:�<]#Z�HB��>_���y"/����m?M�I݉s�W�d�&Z�	EA�1��^�w�[d�w/m:�o'��Jl�G��o ��T�0ub2U�ٌ�6���B�P���Pm��T��H>�����i�`�SB7�"f1��M��,b�U�+�_�\G*Z'K:Sse=�0�S��l��˸V��5:���r���C%�+������hV�iND݆Dw�K��t�C=TU�E�(�!}�8�k��@[M�=��"��"���Z��T�dr���_9̿�C)ƫ	�5�9�����x�����ɻ�gs�%��!`�IN��9 <0x�~����s�oŏuD�Bύ��:����������.%��G��K���E���=]�0�b��FU\M����dj�7�qo�I�46l��z{vVr�m�jBC��؞Í�;��h�y��̔Dv�4��L��x�wc�V����d�0dX��z� �&��s	0��{~w� +]���Ҷ��������Sd���Yԯ�����E�>o­	-���K c�}� xd �V��'L������ŷj5X�������q�yk�TV���7����=K��X�L����p�U�D��P��g�~>��8��M�q���q��?GM�$5'�?��7�?'Qd�s���Γ<!��9����9��q�������~��E�9*"�y4��y^�9��X�o�>F.֭�nӛW�p#~m=�Ճ�5ޭ�m$��ͦ|�fX*�����P
b���Q�E>��)׈7VJ|�O֟5r �R�DY-���ah�6$�V��\�9�^��0X��,!/�� [� �I�nl�t���b	@f�����*m�s
JPP�xOO�xl��@fQ�G �̻Uo9�GrN5"_��P]!�G�,�;xhKU�z0kE���*/�-��]� �Sw�^��������q�����S?���+:	�[Q[���%mL����'ۛ��W7���lp����b�_!��i��H�U_�/�1\pX91�� ��̻�����o�'�ȴ�%[Ͳ�jy\<w*9��i��릦��P��?x����()�����A�A8[��}ۨ�P�=���xf'����.���>f� �0�,�Q&�����3��`�'02z.'�b["	�q7g��&o}�sV�Z�J�JW�Qb�*:��A/�����[K���:��n���vf�sദ��q���m�&yfQ�'��/{"��_ϻQ��#�d�'�.�ʘ;��)I�|�q�8���jG��A�2C�6�xz�Ǭn�/6���Tq��l��~Y,
���`p���s<|Y��4��/��p��Q\_�9�ԠJ��~�:Ҙ"�ԗZW�����\��Rn�M?�j\f�N��@��5�i�w���hw�C\���!���rM����,9��b�>c�S���O	h���m�7tWY�΅��T���0pH��	��b�s�mA���շ�|$K���A}����R.��uK�ʀc0�J����*��
i��t4Eq�� `�4�*����kc�X��T9MM���2��w|�����6���ۨ�4��l�(E|��|�Q�p��w��ab��ˆ[o��*9iͶEg�[u��>3!�'a���T���D}� �����āo�5ޫe��:f3�\H	��?QD�ɸ���Ccկ{��<M������� ��T�n0nBh�"��~	�~gc��Т����}]��NS�C9q�����[����Bڂ�������ӛ����	dS�Nv�c�ĉ�3ZƑ����<�tt�B���f�X��=������������Nb�Y�Flt�J=0�+w��#@�h}ON���I��i�A�.N����x�|�*sT�`�i]M]*�@ᚻaú:�Ƌ赡���ޢ��b���e`��> U1yN1�	QL��}��?���<8@��J.7 ُ�r�hH�P�����H�\�͈́Q��o�xbF/ب�����>��g�=��o�mfM#Y\�n��>� �!�ie��K7�5F�߄�cJ1�K1+����9����xZ���.I$uJO-]�b�ȮȠ��ǘc�!v�3uV��4nJ������'�[Op=Z�Ԋ���(��waD��{����/�W��MN^��jQ]����}5_`���Qf��\�1�}�̼Zc�ևM��s�M5��|��ߢ�B��4�1�{L�4eE:�TT�(r�h^�KQ�0���0���F�m����l�����|z.�m�Kʞl�_��]�_��r�T�.{��H�kq��u���07�b6%�(@(��C��%��kO�R#J�}�;�67��a|���1;���)�#��&�l��6�߽�\1+�$&'{�Q�T?/c��`.�� ��"aM�2�,E��ĸ@4/��(���0��UYcn)/�f�������,�'�&��~~�{ɫ�ǹ����Z���FO�*�����􌾭��[�zs�N[�4u/<��wG$�ߗ81�9`���gh�j�Z"��i*��� �M�ʁg"��\MF�9!�N�HG	 �d�m����Q穡�'�]b������4� ��|����髟���Ft��$��
>��S'��[+�JI$�a�v�����U2���k�����nn~�KU+���I� H���h(y_`vO�� P�ؕ��V�.؄R�5<(1B��@������0��t� f�?�?�݊�r��@?����ZIh\
�$T�h�ߛ��)Q UX���)�E������T�1(���͍#U]�)t������`@$�z32��1k8�c��Gzq�Kߣ�0��b��#���ƹZ�>o9w]ii�F��8$ܞ���<�)q����5)']�y�u=A\7~�t�6[#�,�Q��v���u('A�s+)~�&j�Z@����=̇ޅ�'vtts6�шNC��Z�b�9��zu�G6��|W�f�z�hN��^ڐ�O��e�F�s97�gH%��:�?���Ǌ�i�V�TW�`��"Z�:��c�r�A�v4��,߁~�i�<�-g����lo�x���0��-:ij,��3n���#�/�G1���DPK�� K+������p0���>��a���f���^���/K��yR�
�z�2PLJ7k���2�\�MY�ԧ�1�G50��U�{����4Z���V�M/�;��&V��J��M��gݤ�S�l�t�s�xeL�C�Y>m礴;:�����fͥ3����� d��9}��w�7��坼�b]ыm����y����.V��V�&oϗru&���]��"r�w��=�gR������;���}ȃϬ�~w}��7 [$niOK-�Sբ��4ɻ1zG��]�b��7x�Ž�y��L�����G�����01S4kg���Y��/��q�N���?� 8dx+��^��-�{<���n�����oeaF�6��ۍ�7�����-Ƈ��}|?��\����n�ږ�h�YJ��x��B|$�~�ҵ�uMT��8Bީ�<���57�^yQX!jI5��pIx�j77����_�0�&��FM�XS팧,uC�:;��Lm#=��ބ"fS����s *�@aˠ���w����u_'h1�=q	sDA���� m�k}�_�pÝE�t�#��j601�F&�(I�~. ��g�9���e���z9�8�ٷ@�h'��S�	W�2�ă/e���D�%i^�����o��%K1�����?�b�� ���� Zuy�~�Ƽ>zv�=�'؎��;O������K�u�������]�p̐��z,�ѓ>�	7`Wn��b�ЧML��*���\��'���A/-N��}�	mx��V�6�)�K��ŃEr�&��l&�K���J������~��3fE󘕔x�^zT�E�-�AO�ߓ~FC?^�\R�H�����|UOr���~T�3�h��6�+�jxѽ�U�����@��8�B��6�,��3�Ɵ��v��H��xn'�JB�O�'�Ę��9%�p�����m�����#j����a��I��Q�@�
�t�[�Q��J�B�V`�Tc:i�H�k����Ȋ�Ut�]�6w��fP�6(L%x��"[��.�nxOꙡ��x�L)#z_��J@z�"��o3����y�N|=4����6#�-Y1h���-Ɖ�����S����y�$U��N8Յwd�w�����Wt!��d��7X������85���TrȦ�SC�OFurw�\/���º��j��䐊e@I]w^b�L`�J5:,b{KE�w�5��Ou���=�Ŀ�hױ[��q~)N[H���$��&mD{����'L�ml��>#�-ٝ��T�-s��&�imhV��/q���y6U���P&If�-W��y����1+�c�"��v��͇'o[<�Q�D��j X�n.�ޫ���;j���R�y\�������bo͡i<�㙙�5D�IfUý������_{��g&�8�OܺǱ����8�֣0*�m�1 �<��M6Hn{��mm�h�S�ng���3�M�臚%�MSP�y,��JV���a�kEl�E��R�s�NZ�	,��U�Tr���:e'lЉ��9Q��%
6�r����AuT_>Z��y�SmX+�k�H�#�ٗ'�t�PB��kr���9����MGG����w�f�~�����������g�'��8��x؍'l2�S�ѭ�1N�9q��輮��6���<����N��R�鈴�貨�[$��1<q���If_2�d ��z��l�I_���r�
bw��;|8�^�����m^{�
�MI|譮���tmM==+��� ���J�n]��F�Zy�ƥy@:1Mr����v)���<�ml�D��љM��^��5����B�[}�\#��,��������S�^5L6=�)�
'�ɜ'm*&\1|��ik4&�ְ;s
Us�{�������sM.TN4�?p3���>ps��vm�F�����ܓ���ֻ�X����h�(z���r�q��r?�-h:���u����e�r�h�'{�x��W�b�5bD?x�yvݕ���7����6���r��r�C�w�
} �<
�}��M�3���r{�����~�i���T��D��5�5Y��(�·ר���Ȉ���H��8�V��Ό����"T��Dc�1���2�M\B~�:��Wkir2@���zz� �^Ao���m��D�;�qX2�� ���1U[cw#��;χ��:8C�9Fl[�7t��	�N@��Z� �ߒ��y<c-�l��%��5cR�#�L���'�`��9-���8�	��

A�D�X?�9���o��z"�H��v�Y��;�r1T)����x�s������ϻ¯�c�����3�qF'����֦ㄪ	x����Hp����n�]KTo{�`��h�|Tdj�}"��|6@9;H|����r2���9�F�����5������w�����1�~� 8���~�!�Δ��h��9۽�+rz�������~���Kѽ�G���s,�e�Q@,gݝc˵̯�u0yQ �j)ʺ�mZ��3����Mg�o9����+1����O��C�����H��i쬌�,����Ha�.6i���M����W���Q
��) /']1uC�^�v:�狜����R�6L�/}5��V�걠K̩�`Ô�	�C�|�����fy�6!?��zjV���oe&���އQߋ�G�g�1�@Ϩ��[S�Lʡ�ۑf��p��V��@�b�)�RQ�fY/gn�I�[�^�c]�o��Ɉ@9�"߳^���SQT`�@��͏'-Z\�����Na�&�iV�d�t:�<�X�O���:����z�܎�c�7#e��(��D�Z�7]�^E!�(U%�k�]�����^�2k���L��݂J�~���d�N�&e4߼��e���	d��&z*�,�.;��;���K	�v��T��H� A�_���Y��m~�S����%ߢ\�w1=׫���9[P�0����_F�;�;�¯���V�fsY8hޕK_W�N��iy8����iEl���m#�	cgg`A����"���(߲��[>��~P���$����5Z��x�rDn�:�$�O#pz\�͞�=^�'v"P �,��W�?��Ǵ�o����Ы�xٕd�w���vn�?K��nc,K~�U��9˸���Ǵy��(�
2�W���:a���ɉD���^��k�?�r��Z��A����>�fi�������f�װ%���@.3���հ�[�)����:�>7LX��!�Wy�h����Ф�����WG�܋�� �g��l���|ܿل�I��|��������%���|�e�9��җ[N&�܂�	馻C�<@S�(^�y5�+2Pe/3ԟ�3�"��B��Sˤ&KȞX�cz\_����N>���p�Q��ɞ\sӮd6��6���-�/S
�4�2A~�v�_����*L��{�pT)%r���c �Է_�x(d�����a�لQ����Ozuub�9w���L����,iz=U	��Ͷ��x�B��08
���Ezs�s�����q=|�/�T�� O@��`t�"�y1����x��iqJ��Go�pz#�|��y8F~�JE�X�j��|�S��x{	���M����R�Q�<�f��9p���NS��J:FڻKKo����궏�D<g�{�ތZh�i�����ܐMZ�[�b�bmI����6��q����!7��k��n�߹��Pr����3-NvswX<�V�������V_�~�g�U�r����-��/W��S�`�M%y��}YnL���-��J��Ř93g�����"��89��B�I|�]\���Ʃ:�C|��D=VǍ�T���D�������7�2�j�$���ظ�$�:m��?z��#�.���~�B�gyު�Hh���=`{>��;�w�}��p..�����������i�������G�Q'٢�t�W�Х��>����Ŝ��ϋM�����'cD�'�SI�W&�]��p�f/��������iEw�a�?|��!�i4̞xkg%�2[p�aC�9f!�i��m��`*}��BQȂ�ݸ����
��~�B�e�YCD%�o����={V��E�2C�QuW�y��s�$������ٛX���G��^K=sȟw��⬝�Vf�Qo}Tc�x���ˏޕ��[�ߥ��%�?��~F&�>O��9I��U�HYVo1�Y�z�_|:���'T饕U߱���ϱ�&��|�v!�(/�G鏦IG��ŉ���u��m���zu\�~�{Ѡ��Q���ǯڍ}HBY	�����Q,�N�#6�G��L����C�<�����k�Rͣ� �ȭ��	9��1�r�i�G� ���-63�5�BBiB��ת�5G��^�"	�c�ܸ�~��C�k��.�^��U4�c�A���f���� v�d�(cw�ۢ��v�V��᠑���4O I����r4���2%&��%|*�?�MqΊ|���y8�G�]_`��K�K꿎��w�@�vN���]�Y��R�����hoa���YV?�T=�K�>/$�/Ù��ɔ��v@	�j�Ps�㙙�W_w~��B5!`o�U�����ʆ[�W��l��'>�3�K�D>N������sD��oUi�L,�����a���Kۿf�p�P(�dW�|S���AV4��ŀ�pV���Z��fO����H��E���J�v?m��^0�M6"�"T��*��6��%�$ �H�?�$���h[��,c�(�i8O%)^���͸�gXE��8�v@UGy-�~�V�y���&7�4�-U�����r$c�=�����?n�\)ɗ�<y�G5�ZI��c��[��0g���n�����r�z�H����(I�5��+F6�����fL�{�6��ȥ3;�&���S|9u�n2�Yy[]�y)I��1�F�O�7�o��O�t�&q���_���T��� �m�5֭�t�f��u��ȳ�?J��b��%9����CՋ�#���F��d�O 7z��~��3l&H�%��L,��̈�{^ȿ��s}KZ����һ㏃�c�e�-��&!}�W�'	�[�}I�u�>ú2i�=S��Y��:,my�=-�V�c�d�&��%�BT^����.���<1~@>�0��7�V�S�[`���vQ���.x0��g"B����#�)��
������T?-�*�?w�ut��L�Q�6ʕ'OԾ��|myjg;�vv^!U�h���nr��x��_���է�V�
�����N�o�d�G�e���O���9IdW�+}�rsT���M��q�
�yY^�Y��n�ˏ�ik�_|�-������JZ�z��×x�{���R�E���\%؉7���0�҄%c
�&�Mby��3];��O���XX��_�k�3��C�_�o��Ng��K�/q��d���yDr�r�P�w�MR�{�+���w�y/ݹ}r�O��js}��[�����eޠ+�vB(���Gx&|V^8�dX�T�P'�E�����M�0�Z�
�U¼uN���� �&w���M�$-�{K�z�[��iiߘ��Sr.����{�p�]؅�[ͽ��%1ߊ�ӱ!|��r:3�T������d{c�1�-yY���6��EQ�L�S�(O��h�]e��P	T��׶��ӛ��*�ʾ.+��#�t���`U�����F��[̯�Y`��5$�����~�E�{�ho~ >9�Rs�P� ��X
k�m�����DSv!��~I&�
	?���eܥ��Q���;���ƥk���VĪ;L���!q�������E�gV"Y�>�>\؝�+A7�m��c�(r���N���
7��!���%\.�<(�R����r �A,�*��C<�ϣf2䈙�,gf���r�[�IJ:HnT)Ʌ{��E�D �Ő��27>"X�j�6yYN�y!�@W��Ȗ����#ܕ$�(}�6O��e^�rԞ�z��^�D�c4�:L�t��� \�l]5n5�>E�o�iB�p7^��&��&�u�êby��ѓt�� �ͣW��# �����ȷmM�+jI�Q�(C�>+�lgf���u�f��(*KsR�_^yA}j��;��}}k��u����$jB'r̔�g��|[A�J�9�6�?�؍��*b�.���1���$��$<����2�i�ՒS�d���rN\�Nugi��'[���wށk�S��tzu{ �m���/�k��>�d�\��^��!=�൵�`��'���d��Z]Y�_�Ժ�[o��}5�S��#�)����H��`��8`c*4b��|����1�}{��].��Z���#��퐪��)1��z�?Vױf�K�|D`�K9�V:6��Df��o���}�b��6��5S�ȅ�~�s�Wb�$���q�¨�BSS�����W\����X�;��[��wX�Ωuo���8�a�¬G�;�A����d�v]2��9Ju�)�~�A?�b��S�6+�RqH�5���
��Q�>�
|6Z�Å��
�z���	òq�>"�w��0�p����:O�Q�R�/�ll�nG1\q�c{6�U�&��1���V�%{�q�L��y�5*��&�G��y�,��Z�M���C¾,C����~#�`m�[�C��߃c�[�V��i|k�m���y:�j��v7�i����gI^Je�(	n&,)X6����<�o��Fy�;�$�NNO��΍r>rt5ͩ%�V�T�|��=�4��d���C�{�O�����0�]��O���Aa���8�_���H�Kl������ֆC�_��R"�R\��p@���3=���N���I$S�s'�.����2�/ ����L_�>�1
(6�w�;TH؝�=6}��<'�Ē��rT mj˾F�:��[a�)k�3j_XVM2{ؔ���-{^Ha�LL{�fΖ�Ő ��U##���ѝcr�O�p)��g#�<�=�"d�������{�?�ǹ$^ύ�l��~E�G�����mm�����?#킛�AFePH8r�f�f�-wG��[xM1�̅�x����<!�d�;��%����v�H��麪�	.����C�bD�L�ԧ֋k��b���5g�2;{w�A�
ۚ9yy�&&&'�kk��i���}��P'߼�w馟�O�z}Np}��i {�����AZS����|�SW%�h��x�˗��<����{6:���nsb�5�JvT��Ųq+[a���$�L<��'
�V��W_	mI�oZ���d�\���^�9p�����#��?�I����u�2T�Q}*�!aU���y��������G���/�w�F���a�U���[��_<��6���u�m^>������ޜ�|)�>��Ҥ��Ȍ���_�g1<]K�)�A�����}�Bdy2�GYYY�a�Q
x���������ce��gB���K�����=b	�).��5�z���(�2V3-���s��\���P����ڿuv�k�h��M����q�-)���8��!��a�O� ���ͪ58 m�� ɶ�u=p�4��vnu���~�G|�"�<�?�T@�'!��݈��5SE�S�2�&��K�����Oe��H��/Ï���캹�z�/Z"�4�_����L2NEE�������G~��{o����k�-4ב�a�-,���j�T/�0X�D+�W��O6�=x��[Yt-�
JH�2/5!��٘i��sޖ�aV�`b��O�����K!��d hn��ş�
��%�%�V8D���;��F|N���p����Uc��_�Fy��9	v]5@������m�w���#�N�u�*I?�SܷY�$+H��Þ7(>te:d@�;��x��A��M⼐�T�'�j�r�0�E�.#i�΂���O��)��F��xٞ#�~�N�H�_m�${R%h����^��=���g j�a�a�4�؅��bHc��{�ۧ�f��ك&��� �χFF�ǌi�nc��"��Ӂo&+_�����Ud�G�Pg�c�dg^X��9d0�Z�=Kkg�;�߻|A��Ҩp����'G��@���w��RU�lWU �Aȳ�S���`�;,�X��[7�m4��'���w7=�/
�7iP��5�R1��-O�V����w"Ք��S�nM�?S�K=�?�!-T�*�#�\�S=�wf���^F�9]���|T���k!|Oy�f�����[�暽p�N���[:�\��%3��i�8��$�-)^Jp1)�N��C�����y�=�b� ��6HY(C�z辶�5��}Ն���p��7��0V뎹GN���xn�D��3�^H�٦�m���f��z���.Ei6�}���'"�
AYO��W�p��Ԫ+���������v��K7Kn��*���_�£ׯ�'�L�5��gv���Y�$����P��P���Y}���w�z>�7	�Zm�Ql�n��D������@��m��yQ1$)r�	��iS�m���9� do�f�5��/V����chȊ��w�Ą8��}.����@�������6����-�4�)�eh8�� ����}�'.q|��]em�Y�T��k�5�'-�ؕ=Hf�ȕ�3j�R��_�/g�딾�J6��#I�}�@��d����p�y�K�wq}������j�g1��k����A$b��$��0D��ȈVye�|O�e, ��6ާT(�7�L���������2$2�����W�? �8*n�
}�u�@�%���'��b�����H�j��G<�
�J�������o�D���r��1�z	��x��,�(+ߐ��;�`{����t���a�s����g1�c�+7��;w��WH����ݮ�A���A��𮡜�h�[0��		x>�5�f��v�K�D���~�g���d kw�o�
�Y��wܬ���m�}Z�)���+-�X۴i�>��G�z�/'5$��E�v{>m�[r��j8�*6ۓ�M>z),pteZSgw�z��˵�%O�{� p�R���į4ֶn��d�'�v��������I��dݛBYP���-9t+�K��~X>dV �6� �1������Eڐ��Q�/�/��hia���EuFs�6�ttt\/(��@�5�/~�E�sA�d%�B�^j`pp���6�P�����Az�래a�> l�V��	�um���/�k�>u/_�UK��YL�	���H�m�5^�Q��7��q����K�S�$�ϝ-H��M������N�ǙE�k�7"�u����ȕ뎓����J�
\�9�x�E0s�5���UQV�m���ꕳ�Gm�#(
�-I��A��o��eݬT��a<z��1����%o���p��sh�w ���6t�{FF��G����$��i����w�ES[�5�{�b�:��;E
��V�����-�J��G���y�`�I^,i*� �� 2���3T\��Dy����OX>���eH���A����[J�`="`:s��)��q+��r��,���Q�W���i|P8�0՝;�#l����-.�N�u\���'��ld	4����եߋ�s+h��x�ro"b�}�e���@������Z�Nc"oJ���A�7��_�����0���[���1���_L!/��Y�MGH�	��䛳� ��Q"��vdo�{�h����$u�Q�@.|_x%��W�q�{w�qN�I~�hM�1����O���d2�r����C����A��M���Jb[41~:F�T���R�i$�Td�����=(�`)��{�
��G����\�]T�:@�����r��^����aPY�LͲ�c�އ�����<�}<<t*xQC����#�!���r<:\Rc��;W,*����X?X�x���<�Pc%.�r�]�F�;^�.�Ǒx��b=}77]�U�y���
n������'�Ӱ�wx�R'؟؋�h���vc�f��Q<����	!fn4`c5̑�$��ʳ��id�$Wɖz��^m]�p(w�GX�\\@�1��b��k�7��MuB�hZ��_qcأ����e��>Qm�DiL�������f��L���=UL �N|�4RgV�������`�8���Ʈ�K+��/y_��7޷{�A՚�����e�:'Eg�ϑ)��"��S��>�tYt`x�"0j�!?-�����V����@�HǄ��x�s�S�ٽH�����4�#2��m��:��j$�J��L��L�oݽ�����"�v��� O+�Դ��My�ɦ���|\�v���q��b�x"��FtW���nA<�7�4��^��]�N�ߨ�(�Ҵ�I��������wn�̧6i�i�pu�.��M�V��I`P�08��H��>�(2+|>��=���;��7��n���N��8[��,�:��ੲ�M����2�6W�g�X�j� ܬ�C���Z�b�s�ъ!��g{ko�����";$r�?�f ~��\�6�u*�JSSS�ƞqbr�İŧ �j�<=BT��U�thb��N���ņN�#�����GL
?ˋ����t�W=/�:n���Ȫ B(7����7���a_�W��&�06�c�p,Ҫ�Za���v��oF}���
�Lqw���)�:2�QZ��9:6�_[[{�`L�~1�,�K?�tw��&AymdB�cfd��R�S���pݦgN�?�x7��P�~�Ɓ+d?�ɥf�|ڂU�}1����SY����5���턦�������W��f�F�jFx����!����tL�G��W�*�PavB�Ѿ�{�U�g��d�(���Svf��n*����뽫ч���F�-O�ǆ! KtKt�n��/M�/�~կ\��#�<����y9��n�f�~��M_�P�η��~oL\ϸ�߫?ݪ�f��v������%��	�d#��I�ɛ��1!MV6�>�Iyԙ�8n蔼�VdV��
$^5��G��������n:!jp������+�r���'��I|����RK�O)�2��>[�4ҼE/���)W�/���}���2�L��
¢
x����]O��8�Pm��Ɏ�\�J��P�8R��S��bp��Kx�^�=^S���6���?j2[�D��Y�eˑ����Q%��_�����g�'��y@)1������6
��xT�x��ݱ~�D/�	��KjW�Rzܻ$��J���j���(�yg$c�n;��Bf��'��1���s�ͦe-��T���8׽�S��������H�gc���5��I_S	a�K<���e(���T�"�{�=?8?�k��G�Ee��,�rI
f�lm��Q�d�;��~���+F���ƪ�Z5|]�N+.��2\A��e|K;�K� w�r.���C��<�a?~SHI�W�Sp}$�J/����p.u�,C�fW*Z;i�(�{���p��ȳ�-K�&��� .��)[>==�FH�u�h%"c��$����y����-yړ�-�@[�k���=�oiy��sf������y�-�z�=:~��:㱧\,JN��;�/�WQQ�sz��CЦ���`��3����{����#Ň>L�{�f<y���_q�����3�x)O��[<I@�D}�z_�4��w����;���[H}�U�.�ۼP�}5e��wjX��&�1#+,DG���ڄK�d��2�ζx�1L��%]����������q����z~�a�R�1;���}��ϩh�Df?}n�����Q':�v��R��)"��p.�q1i�	ͩ��b�J���&N���D	�M![�����~���L�t���a\pZ�h������{���D���!x"�+Ap�(�pY�<�e���<y�dd����9�	�l7���=4U�e@h����#��w��DSs���df^qژE;��YY}��r���u_IL���a�g}q�E���#R%������}8�F�g��|�W����4�ЁbU^̜azf��X��苷Dw���OE�ʏPG�����#�'�v���O�����e�v�2w�����G�ҫ�t����Y�Tf�:MY(uq�<jr�tG��$΂�}��he���f�\��v.�+eK��Ǎ��Tu�G�Q�Oyq�fIC�(�L��x�o,���)��x RA�ٷ���RU��$�^�Hr� pD,���}�%�[�(0w�+p��,f��3^pӪm��E��^M����J]���ݏ�w�Z�ͫo���)C�ٵ
0u�����]�4���~>��A><<<Vb��p�Ly˄��|�t8 ��ՑlG�Rin0������)%�uB-(���ב���#���t��Ru�|���+L�1;��h�ӪaCRg����뫴^����wno2�P�V���MI��k���8�q�"�N��u��sb��bp�}4������yv�}L�$�[��'��O5o.��z��R���65RhYӒѮ|���~2"�o�\h�_>P�_���i[���2�p�\��@��b "�MJ�� ��jU��s��P	�(Y�ʏ�M�)��)���]{1����ڹ��J.M;�7o�c_�X�`_'����Pޛ�&�u񥮎*==ݟ��R�hz}�m@Q0EUWW����/P3�s�p\^��Y[�Y��A��Q
2&H��� (T-�)+9ާ�TB�����SQ��j��~33�G�������1�,����;l��ᛓ�ׇB�~�Ҩ�͗�+�WP��y/��v����Y#�5�.���Ol��Ll�ҡ;B�,2G��܆C�%�0��f���6������S�	/�;CY89Sm���>+�T���'q]R'r�R�$�o�}��[",�s��� }�����U��;���w^�E,p��HuHF�ܲ��+ϸ赁�F�ߢ����<pJ���m�83)��l�9C�]��Y�L�@[I`R�w�uk'��pe��z�E�ϭ��Qb�~+[z_9�癭�?������>���"!�"H��J���-!�ҍHwKH�t��đ.��Н����{���ُ�zԳb�9�kͽ��ח�!����V����&��}�v8T��Rr[/ϴ��f �������]>k�mAro�@Y��IO�f|�L��x�c����s��\��č����Ɲޙ������
��L�oW�{'���2an��ܝ^��XQ����@��ի�I�0=�$hu|qe��
GFN����>��Ņ;;;[�T�=>s�H���7w���P93yId�AB.��9&�_G(�3P�!!X�dX_�*��|s8T���W�N6$<��L��������4�@��N�=NW~�𹽿�Ә��X{#���'�����͟d%��~��	[���R)2/�P֎�Uib��ob
9z�Aٹ���\k���;9���8���׍Π�����n�`���&=���O!��v.�U^ẫm�!v�w�Ls�q��,l����FM�1�w ���@Q2yab5�oo�iݔMRI�r�}�3��'�f%�U�'&N���u- C���3���<�XJ�ڵr��;1����굧�Ѕ�>t}�������퇯#K��P��@�F��Kh�dߥ0���fs��Oɥ#�5*�f%�L�Ϙ&�|�����y��_�F�#��݀������e._H4�Qt���
~~�N�v���?��#��%�w���g�%$)u��3%.Җ���@�>�2�@��ǀdIBBB)e�{��~��e�-�-%-�ee�J�&�%5ޒQ�&R�>0�����ru��_\^�Dw8���h́��>��\�z��U�"�oL�ޘ(����s��&"m�F�v�/LZa/輏"L��ƆzB���11�
�O�ϥޢ�ƚ8y��H�|u�r8d�Z{F�������ؼg���'�S�[�J���m�ɷi:�<z����wJ�@̱���$�v�����u0g�wg�(���d�Eȋ�(CF|�<��Ȝ#pK�.�?�[������(뭟��Ò�b;��I��8�4��YC`� �F��� y�椻or<�LyĶ������X�H<A9�B,	�b��of��߽ٮ����{�E�d�[���վ�����s�׷{�>� E�Nm5ʞ�b����X�`��U=2��J��o�gd_~��}T�k�B�y	�H��R��Q/jy�Szv�G�_�P��"l��cض���/�{#@�e�E
� �{�>M��[��v�`<# 䖺����[l�@s����he}����P�f�7QCwߟr=8މ�{�p�S���;����+�Y�o���F8"������F}w��3��(�I����H��S���MR�-�,Y�P�h<}�ڮ3����8��}>�s��xG���Pkzz쌡Ȉ�����|�t���������n�CE_D|�ˠ��0�HE�u����$�>z2RJ4��bX���jd[����ǝ{�=wC'�����JlP���AZ}W�����E�i�ǔ�B��ժ��� 5�J�6i̓�b�,w�W��.k�><�U�pj���7�B<R�ጿ) DMMMw�����Hd@ɗ�`[�P�[|bo���g��F�?� ��`�������FZPwD�}��m�pm��WzǄ����DPP�߻w-�����1���>�
���Ύ�q�5x��֣��D����"ы�i������p'��s�a��#��,~�P���f������)�%H�5)���ޮ�ܨ˜\UE�H��>j�޺��>>M7���rX/j�d��e��7�x=.�V߆��J�7O�A"�޶����tqqQj'�4�� <�2)����Ν;l���,�&��x��tyKC��0������]�?\�8̌��r>F4�Ӭ-�H�Y>Ackkk���5x$�j`]�X�M{b0|""Q��`@)����00R�����ݿu�Z�/T�b�aaZ��W�y������Y�=W�[0�v�lSz�_�ZL�].F���1j��0H'��::���T�����d��������Z%/�?�\���e�৑�U��U���9���B�f9��}K��?Q���c>��z�����p����7��@�Q*۸��(��������B����A-=}}�@s�@�P]=��X��oy���9S:�1�ߢ�ˀ�l1���Xd����x " �/}: 聓����B|G''�хg�dd��Id>c��]�����j�L����k��.�iK܄Y�Ӡ�ِQ)��o�����m!w��wD��rpPj��f��P$�3R߽	xRz��H1k4�ߠ.�h>!�'��P�e���:�]��M��5�;�o������.�A)�^	C�6�����<ߔ��W�iyG��=�=S4�3เ�n�ˑ��G�0���XqG�VF��R6,��G�.��X��0;����Բ���i���f��7`�u�M˜������[��)�g��xcĴ��`�A�o{j++	&��7�}i7y���(�q��$N�!�RPP�n��D]D �ϽD���"51����C�bbbr����f;�ԯ���*V��.�	�����X��������r25��;hfL���v1����i,����Y9��8�O���0Hw��_�� ''װ��8�������f���"`����t*%wy�z�6֪�g
[H�66,�yn�0��a�^�i�FA��|tt4�i/b��>��|��w
��jA��,��>����)����1!ǃ؋�����|�*(���}�ؼ~�ĕ�K�ϳM��^�Ǒ��0qOL�O�w'���&����w?� D�T���%9��-�F��G >����߃��0_�b���� �gb�c��.�7H�1`500x-.�����+k�xu��U����{����ρ5���'����Q
?�咈�J�NG�ﱿ@�~Y��@WqYb*=a"~sũ�Yy��w�:� ���&�8@������c�7c9�T �ѽ�{(*'��<�Rw�g!'����uy�(���ej��^l�������5gG+��$����^B	��s��)����\-��e,�������Q��uH�����@�c:��`aQ�!�|<���>���e�s��)�T��Jnl���h���񝬬����yZ�9 !�YY�>p����������@��@�zUK�p_^^�ַ4eUiф�j���/>L�����7��c~�yI͢���?0%� _�8j��z������`���;H�\���DX=b�X	;>���<���; �f~�&ce8?�Z|�Xcy�e������>y�Qq0�o9b������l�d����V��QdH21�`Ee + �h@�� ��IZw_8:u��<_R�4a��M��Ұ��m2R����uQgA�z�&�ņc- n����W��Џ��U��{r�e��S�c�!��X=�k�Oo����|ҶQ��/��*u����ycu��(j.����B�����AxC���1y	Ւ���M>����_G���i&0<�����C#���Nŗ3�=^e�Tj���tݍ���b���$2������x��
�<��
2-�*���lox��z�(5'5D�V(��V��֗��EG�W1����m��Дs&H�Y6��)]��G)��g�?�J�'������6v�!h$�̼</06�u��	v�H�\݆���"CM�|�Y}�.C͟*�k�2M�Z(4��4/0PO�W���
ƎQ?6��<`PdT��A�4�>U/�����:,���v��1��7s�=���~(&��활*,,��#��M��_.%T��R���Cו�"wk���p�~�@s
�l�H��� �W��m3eu�.���)!�F�N�ޱʑO�=Z�4�[R>�X�_��5��tDZ9��,����ga;�� ӗ�}�9;'N�K4?����OǇ& ��1BĞ�t��xzz������r�h�.T,$:113��u�~+	~a]�+�6\W�τ��?���.��~@ $���ڍ�Sd��J�,Y&r�Rڰn���ŵ`#�'%����������(5	�J�^�F�Je&k��cn��ǈry!ɫWB��ˆ^�%qv/�{��A�&d���Q0�8��= t��Nw��(�mm��)X�;FE�YyjY�K�/�)K ,%�I�>(ۇ�Q��de=��U�S8Y�?�U�S�:^�?������W-p����z���>c��Qxz0�.w��^�4vU&����H��	�����{=`&��ʣ""�KKq�ѕc�y4j���	�(1�Hf��vO7�~��َ9��*UZ�=�}p��`ra���������]�i�_1F��i �-m�I�</YY?766�"#9e���7,Y��<���P��38��(&�����P���M��M���6�k��s��}@������%�eC��αo��Y1g�������:�
:��
�n�F�j,Q������ E���$Q2��azs_J^��B)o0w��b��}W"�����Ì��*Ԏ����W�z��	
��h�#-�9.�>��م���l�q
m*c�+y` �a�<����V$| �`}��MF.3��`(�7`�n�bs����.Ƕ���� ��Om)���z��Y�K�&���4�O.��txr��eP�t�1@�6f�')!��(� p!��B�Pʷ��)|?FLq�^�������bl�a�U�6ݟzQ���xӉNk�St�/A�	?ොq�g�?�5������k���G���5 h�a(�izF>�>g���>8��?0P8&!�  !!a�ؘsC���_�D�����Ȱ\�R`���	����-���U�V�(j
��|c1��9��m��{a<85g�ݷ���OL�+_���N�[7 ى~eN��C1���н�?`p����G���p��M�H=�¦U͛��E��~��C���� �e������5K�X>�U��C:�G� / 5b�ajJk�U��2EEE}��b�͢�=��ꠊ�J P@ ���qC��!��Q����b���n��p(s��bN��멙l�WD�(=rt��Y�^��V�]��s��w=�/��� 芑�?����IW�h�_��	&��}���{�S`����Ot�⺇.�tѻ,�w^V��EY��<�;F�L ����#���;�;��֏C�t�sz.��YY-�8{Р5��nw���k�Aƥ*5۝���sQ7`����7��K�o�Q\A�2�
�~���{��-1B���F|Y���S;��~�C�_?J�yt�Hq
j�S<5س�&��_����{���Ǌ�O����ȅ�JJ�g>�����Jr�
��V�Y�S �AG�y�ݽ	�w�N��'T��f��cu��$��Ey�+/,� ����OK����(Pݕ�+o��d9�DTD���uS>����I{�Iz"��H�&�TҒY(���d8�*�\�"yjNz��-"\�sk�9��E8:�O��E�`�s|���ԅ	V�NY����,�m��?cK�`�QX�ڒUu-�Iܿ(w
`���}3�g6�^��}��U�	��h�^L{1�xף%�7^�yV~\�iD~���6$|�fT�����J���}�[�y�5�� ��O�f�-�%a�wv%T�Bf�_U�I�j���Ė���a�����
A���~XU7k7����ZW���� @W�#�x� ^�S�`	�z�>))�(Hk����ӧ�� ����L�핿/TB!���0��H�L4d6��	��i �V5��<�Zq@�%G3����xϰ�r��9x\f6��ȕ��W�ߣ4n-aU�r��+�}��q3ff�o��n���j7�����4f;j
&՝������o�O��UU~���A�E��c��˿�/+9�i��'�#����ӗ. ȗF��O�+)��_�V(���=��-/O��E�y����UT�Ć#Z�?���~`#� ����(x5�F3?�xBvp��@� 8�x�xV�� �#*@0!���d
Y�P���*�<�SU��4�̗�D�hR�U��W���v������g,��;�K�#Z�d��s�Y���^:r�{O���^�/Ŭ��9U�HX=y-�}�q�Ipt��m��u��rJ�K�xq©B�ʐ�/�:�r[��f,;���TtYvJ���	D���f�ܮ#���΢���-s��F��no�b��b�y�ʺ8y�����g5�b����jdb޵Ї-ɕ,��=��ő�4�e���Ԝc����/\�NM�׎�~�Xw���?N�Ǌ��e����@j�t�Ç9��"�A-i��Ɔ�D�#C��:��ĖٞHz��u�����ݜ��b$��F^?#|Ѩ��Ja%����)��#���uU*�YŹ�<� ��@Ǖ]Y^�	jyG��iϤ#�[��=�kB�gaGs�z�2������������ǯC����pͳ"����˓ob���k�p�� ���')�_��������\8c�Zh��p�;i�@.� �����V��`�&�k��1�8hw��ƥg���n�ӆ�1�n�;�y�϶:���� ̭J�c��_C��@pyκ�_k�U�(bp�t|r��F��f�6///5p��9�׭���X�뵷��I�ۉ����W�Wh|�b9n6?���p̪;E�����}�/{��UޢK�L&��&r/�I��B�tw1�r�Z�u��>��T�ecc�@�_��˪�R��c67/p�
K�,+��U��(�⡅�|� <=�<�u�I����S�_�M���D�"W5]^�
k��Q0���i4������>�劙my��9+�r���	�:N{=,�'�4m�$�{Z2�Y<&}���X�������cƋ��ݳ�n����0?�|<y^ɨ� ���mbbB�E<�G�X�+�=>��6:x/mAMʐ��i?y)?Y2�I=r�I.e�B���lIN��Ą 0�ʥ��/�^@�߾���-�pn����t
��;E�_W9��@4��71�IK'/�ep�?h���cq.JS�9������.*Þ�#�d���V\���6d.���si��ۆa�R����c���jf����-��"��#PPQID�ie�A�S�lU��W�D}�����i<���kg�/ق��(��/�*�=s��ڮ�������B�"s���z�M��/:��ggS���m	Z��=]�|5����J�Er��2���>�u�S���ٍ¹H�����7+�\Ը-�B����j����˖rr���a�,.vK����� ��=?���, �z)+#qF��-6�2� ��8��-��>W^e]�=��h�b��w]�,�w�-}�8V�q������v+*
���>I�<��X+��������d_X��L��6�hf
G9�����ŉH2>W�E�w�\�sC���
وI-�� b�+ ���"x*+��9jftMT�Va���4>���tc�g�kW�V>��
��ֲF���C�(d<�a:jd` ńOl)fk[���)����D�=�/^(���vq�ǃ�x�+���}A^���ҥ�ei
;E��"�|K*�)��˻^�����R�zjQ�baa����,���o�܅i�����]\N��41�}�&0���Zɯ&n�t�^8��Ө������u�!H��cV��5["�ey�����о��?>�}e����w��T�/��'�C��-�rG���O�Zf�ΎVl �c�<:^$�w�X%7�l���y�k`�R���]O��1RZ5�J.�(QaRTTF{�H̳�����څ���^�ac���ngʑ�A�P%zib���qP���ά�Ĥ�~�%��R�N��?0���=�>ZLeF��@$IaR\\ �2f����	�Ň��AC�M�P�5�k��ui�iFԵ�����.����٧1JfI�Ne��3�*��J��s���~��ھ��VDY������O�H����Y9`����u%_���UTLg�{>#*��"�o\^L�t:1)�`$ @
���:9qI�� ��1����H�Pk�aSJ|U276�[)��_]5��헥������e(���ة����x���E+]@W����VT��0��E�3 Q7 ����1(n�o��QVj��/G�=@�&���}�/l�����6�Om�T[�țZ�W,� |
D/��7�J�k6��X�_� Hs�{�YF�%�o�����W�f��)8����r�^�� a�T��4ŕ�
¡�6�G���
W�Uۀ�D"�x�9+�,��)|�nUc���?,���4X�eU��䝜�
4�8�k����|����#xv����%0b_��І��y�j"����4
�L���RVV�xv���ӷ�$7�i{���
�N؈w�4Љ^�E_F�����e���m�Ћ6Z��7�F
rs�=1y��Փ��!�`A�����r��hFr_���nU퓘���{^�Vwl�0֔���426&�@��)y�3퇚2��vL>\��d��bBbs:,*Pƽ��������V���7�ǖ�B���E3������R=ǥ��_�ж~����!��m�Z�Ҳ2#--�_g������ �:3
�
�N�Ow5�Kњ�YY}��GfUK�\�G'�q������݌5Q�%?Yj�NC�@���*�񔍌����"�e�,��T��2�8D�K���w�ხv��㸼�f���=@d������:f��G���d�%X�22qwNA�v^A�$dwCì��u4I�K���[o��hH�ք���§`�\(���t�A�ոu�(B�)���XN���4���`b���Cȏ���G��H8mŠ���S�ת���N%Sh�ԯ���~�ӣ�޼��ap�I=�&sA�"���ĵ�CG�,��u�z2��)<�PV�]��IWU0�n�tS=�1���&m�.�E���U��������
��D3��t��HS
]��"�M���2=t�2�a�_���/����f�ꉳK�7[ld���;�ϖ��V_���5iv��Ә��x\��]NW4�c�$J�G4�^N��nl9�
@n�� �oĹ�5u�3�e:�U���=��k��w�B�2[���UnT��UpL�[���6��,�H署o檽��3N�ܠv��$���b�
��"т�9E�Gi�f�:��x��,$+�F�mk�Ҿ��WB=%�s����(x����[Ps������F�.3W���u������A͛i`�-S��4v���ȯ�V�ꡕh�"ٵ��F59�����]Xz�=W���VT�z�qxT�$�> ���^��7�v�\�bgU/��I�p?=�"��ʛ_r��n>8�$`�l����ez��O����?�&AH�7���0��vg��k(�j((G�U
H��+>bA �VP �9�}����f������u#I<�	��g@gdt�gH�ONO�;i"�M�B44�E�*��q�[YXH����f �<?*8_���0~���-@>
g�)R=��:���}(���	 -k��'b(W�P��WӨ3�ݘ��*bO�O�]�J���U3~�@åm>�����i)��.x$}մ79�x,��b�|G\m~���=D��y��UW ��1�����3̑���(���S�L�����
�R��QK�p���G%.:�5��	������B[��̤*�w���[��u<?��1�Vc��1��';�K�4B��YLYÑ��7���p�Fr,�]�	���[+��*0��ԫ��頼BH�z�쨪+pS�)���O��Jz�s!̓}He@�TTUA��޷��b�8/��w���p�MN )7��(���b��xu���zg�:��[�]��b;��E�#����遡�����m:Z���xǌ;Wj�T�s�g_�"!Y�����	�p[�Nގ��e�<�Z���kk���\ ��њ,�H`i��E;+��*...MƍZ��sl2n�'��~}?[G�;�G�Ri�?ފ;�*0s���������<%��,W��4�Y�Z�-x<�ŵl� �UmwrF����2ט�{���y�20PH3YJ��d��)9��7�B""�>�W�,à�>�?-4�+��d���W�>��x�.��u�W�Ѳɮ`��fc��4j�����%�4�;����N���(��Fff
\��&h�&����*@~�T���h'�%����o�bl�2dݩB�y?���͚Jd������&�8��s���^eR��j~��Ū�*V�Ek4��2��٣�`����,PV1. (��k���R�����Fp��ڿ.3�$Au�]�iK�<���w�<,A��U���Q��"����_�����5@R�p�3A��z�a.B�x�ݹ:'G�x}�a��mzͺ�F�ko����Q���M?��@�%����N���d a�j'�pIL�w��B�H=a�X5i�'}��`L��w�h����5�t=6�z��{��B��+1aS��
2������ō�n�~���|ౖ��F�A��]��{1)�}�+y��55jyyy h�V@���{�����WPw��a�Ǻ�g�������v�,�	8�
I�ɊYh�v�{��~�8�\�
��$�PS�Q����{�@��W�޾y�������5"2�2���xu�����(p[�� *u>�|ՖHiT#ΙcC�FE8H�a�����d2fj)N��ܸ���V�;S����%%_��X�A���:�]S��@3ն�����0�ɓ����C�5Pj���ސ���w�sܣ֥���-�_]7M^��z�3�R���ۙ3�-��]�ܪ�A-��L6���מl���+� W��ӫ:��#��><�@�"�����w�eM�fLh��5�� 4�/	5�]����$�W���d!_889}����奤�@ǣE�=;^ǜĸ�9Rj�_��:�?�9	ss�h;�Zb��]�}[����G���������i�{C*P�����2�MK0-���Gg���ʦG�}Y	�0���[�j��ϔw�T��0i�S]̤��(� ����m��b�5?/`�M��98�'�-��3w4��G��, s�mK;;�<Woӕ	��7y"��Gם.G����ʒu��PZ�%�(�7�fD:ChK�0�����������Q�nګ!����߿���Y2���剛ן�m &&4Hح�E����#�*d�qQ��f�Sv�@2f���RN���A:��Z��˩xy5��.�M��XQ\6��P��Oh���{�����q��+�s���v�v�J�͠{���q�"��J0� $����9::����i��fP���D���dZ���Z���z��#�ZE���U��+d{���b-�r�0�C�1����r�>K�{�P/Z��Z��� �N�L[
���+��ؙ��j܄�1bz}yy�W�nw"�:o���o�#_�*a�<mM,v��@*�@���[�gK�K��T�`7�Rj!ϖ̯���Ԓ��e�����ި���L3=}�a�#�t��Q�Rg����5�U{����MH-�ġ�okEn���&X�%�e!�������ْ�ВF�2�Qt�Q�	�"D��)��hB^�t�3ri>�G0�dXx���>/E��[��/���!�#bI����**�+��\�D5e��d����،��b��I�Y��2�kU+`-�rO��W:9����k3���Y_�u�zWY�XW�SD��;�{�x2%����V^q�r�7��#�(pqp2�r�q���J��,���-@����AsQ��-�fލݽ�,���os=�"��H�ϰoEv����xS:�ϴu���N��Z�#�s�	]��OQڀ���"Q�-�c�I�ÓӺ0w����o@
-$:�/����g@�����]��?�����T�}[�[b���ʶXy���F`Y1K*f2O�E?{���?%�g�BXׂ���%���h������v��q�r�>�TC�W����z���Ԁ���JM�:0s�d��f�n`�s�ׄT�d�LLֆQ��1,��h0���ɕ��N�����8�� ��7Z8��͑IC�n4d�����ȗd	:�|�C7�,q�g�Tp8e����"  @CC���]�g�.cl�H�$��p1�<�m�Ɋo��W��Y;���P&m�[��><���.��:#E�U#^��H�k��-�'� ��b��VO�Ji�Ւ/-��r��l�:l8���f��iV�o!*þL{\\���-(�.����a����Q��ꥆ��%�=L74� ��q$��
~�t�y��蹜蟂�1�9�����T�SU?�W4k��%"4?�4O�.0�+3��c����~���i��&�l��i�P^.~G���!��~0��Dfo�7�'WUqd�^%�׿7�E���
���A�g��֣*A�%����h:��^�Z��0J�uI�!j̬<\�Ack�U˚�et��z蓌1b�EP S<��z(��X:���r"h��ړG���r�����j�V�wxH���[���xw�v���D����V| R<�`K�4��^^\�� \5i'��-�׽��3��vE��t�d���dε
>I���+<N���k�Y4����VH�E�O�c�!����Zr�{��RM��h]vvv��"���D��+(D�h�}t��ԣ��� ��hn�����Փ\]���sJCMF{R�KWƣ�vFp/8>T{\ٻ�<h˜o���%P��:z͚x�%�r��=�v�N����H6?�a ����4e~:T�? [}j��pّb�����}�O����e�*���n��7��?y{��hX���i[�YmYʕ�*�2-�''!x�z����vo�֞�sqY�$I�$�?���YZL�RTi��׏��~̤�qB�����n�����$Y���uԋ�m�F㎖��{�*��ü�	L��*�?+� 77w�w"],����,@�g:^M��R�������|0W�F��t���Y��*�%#��#."St�ۃ������:S��K���\8�����5�������k��67<g��pm:�rǓ��Z8::��o�X�h �h��T��T���ռP���c�ex�}_������H�����wnh]]��� -���P%DOO_d�*��BD��X�� P`>�|��� �=��B���wFaZ��n����_�Z#S��J�_��ț��5������{���خ��f�^^^4tt��=iO���3:���D	�j

�fgiU�zu�4j��2* �8~t��"A��L��Zہ�����~�l��K\�V( ��i�b�}��c���`Fȅ��R��q��G��v�f��og�/B�Y�Ӿ�w���\e��F���`V���Ȓ����s�[\J�im��b�(���礥�SPP���������@7� ui:J��/egW��f]ee�ȏ3f�`��n�������Y[Q�ӝ"-� Vm���`r��<�˥u�PhvN�M�퇙YY��l:��bҗ,�a�?�DU��L�ǟ	�T~� �5O�T��n� �)��:�w=��٭`����֥�-b�l�|�}��)quyaa_++���U,h|�o_�v ��&��40<|���/��)sh�z�����E�?M���Cj7G�Q��ja[��ܙ�^ǏH����ŝ�p{��tS�hqq����?0ǝ�@���e#a��%6�|u1˫$�n���k+B������DO���q}��x�uK�4��6"�ێ�Pו�c�>~�<>� �?ߙ ���ܿ�	�ד��5kS�J���rҢ�������Y�^���;�E�2�'���֭����Q�q5���/�v�`wy��ĄX#���/���2�����2�V)Ě���/����¤�:_��#^�7Ş�6+����:�g���ǆ5_��z��"HX�i�|O�����n\�_Y�}��g�f^�-��B1�7���v�%��H7��|r�yLY����&_7��l��}v�*,���#K{�WZZjğJ�s% e��ֳ�d��w�7�����7��YlO�e��X"��E�䭭.�eg����	X>��n�Ꞅ�ǧ���~�ғ922��ݞ�g~��ʐz�?��Y�#CI�X��1��������p��&���׀>{_m"Q����^�-(f��	L+�v�7�J�}!ȼFFF���+��]����	������4?WII��y�3�rw�Y�ةli��LDO/鼿e��""��z��ٞ���r���� FB�$��n{6>�=t�r��ü����L�8ρ���Cۋ�	g-
m�r�Ȃ��$ ݄C�.�{q~��@�4:�a�DbX�,������C�	���IÅ:>f5��>�פ���a{�^t��r$�	�7�o��E��	�.˯�����p9��>��,X���$|W!_-�hT��oSi-���˿s
���3�烼F�+�b�˫�j!�>�-�HY�WU&?~�|��Z.�Kc�,��>��pXH��������24�F��X�RI�sI<�U��Ŝ��B}�:�����\{��j1p�W��4(���&����uj��͔�� 5����Y�E�&�4{:�pҹ^�Eȥ�)(�OY�_��Ž45�����o�r��B�v��a������!�u��1[M���:����?�q�=�Ӭ���uc)�##"��!�� ��A2'� �~��rJJ���xtJ�ޙ���0O�=j��%���f%)x'!�u�U礁R��j��Gm�(�(f��5�4+a9�o!�CM�B�����{�G�(��k�����9 R%M޿O��w1����[[[%�K2��Ur��nt@@V�D-{���ή�r�q7S�� �[F��ƻ�1j�Fook���LJK�l��Y8(^�-�������d��fN�ن��YT����"vA���q�n��v�/��q���cP��\HI!s9,#*�QMmX9�յ�L-�6Z�{���,����'@��տ���)GR41�)(�[��ܑ&�ֹA8 �I����`����e3e]���R��v'*Ǥ��$����R�
m�;���```@�P����/���%��t�õ�J�B������C�
mN�R?��q(��G�pyih�8P�_ժ��S.d���8-y	va=jC�cBӄ�S e�����S�А7�;p��&" ۃ����w�p:W����3���I���8�c��hH�������Ud��w4�o
��v������yA^�}�Uo��>8:9A���/��	c[�ݟ�%	�j%��z@^qs��*���Bӑ�_"6u��� �j���V	��p�J�`�E x�c����������5?\Ǎ����3L�Ra˟��m���\B�מ��� bW)�����"��$j�9��C�����Ы�������tUʳ���F�
���TJ�?sV���TJ�Q�%�`�U����� �wJ9ͺ��4��
d��L �p,=�V�'�$P�p��"�@��HK�u��܃��0>�O$��bqz��W-j��)����{��t�t�_��YG9�՝�����/r�I98T�/M5z��(7U-T�1�>(6!ДDp���Ǫ˷���Eڵ�3�P�A��c��?݆���iYHH_zS7.�rK����c+F'%o����\{����vM*��m'�6�+3?~�Ḵ��|�.�G�1���-7x As���l�^��]Q����;h�-�Ɖk= ��`�L�o�--�UK���Pr�fWw=����5�gU�=�4��#��f��p��r����Q6jI�����!݊~颢�ۇ�	OH�S�h_���N�r�I@j0R��?ȧ�w��/I�x6ٮ����-��g�ߦ�@��1I6��*���,oo:�ܺyq4)�Ҹ�� �:@��L]�z�X{0�/�r�bL ]��'~�� ��5fS�[B�x��t��`KZ�l�el����I4�S���(Y���[���*BB-��B�B�	U�9h��������7���8�I~d���15Ed��jh$�Vl���Ffȏk�yE��[��3��(7�tx��Δ��	1$gv�ڻ��� a645�wq����-�[�P�l�u\���y)��؛�p�ފ�n�d���0(�v��	*��X/ I�j`8 ���Ը�yÀ�𸱻��UP 	�Uf����o�R">��Йgna!'3SH@@`˞#�ĺ/]<lr}h�ɧ�n��F��8��qzW͢������^E�6Ə������bl����M����Ms�7`Y���/��!hg�S*|[m�nˁ!���D�[ng�DF*��+-i��e���y�p�e�8��k=���5K����P����(6����Ձ[�@��2�$��O` �0්���~���4,XT�m:����@�cc\Fn��
�I�g���MC}��5�飴�:���;48�����ᷫ����{0�{$�B������	�xIl-~��Ƃ��	<���hg5����j�U�M�I��瀯mE�綷�w�����A�U��v��9Z���]^]�377��~|_
<�� ��̟�x;��w2T����SV�Цk��H�:�o���y��-ؑg���ْF�ϓ�����=�Z��jU�E���qza@�C�sP�bh��<�9G!/������|�ɒI��>��R|a�/�ƿeI��$���(y?V�� �ѝ���3���P	��#III���sVByQQ(l?.H�x���4���8B~@�x&���'�Y��<��)g6�bJ���3����]�����l���޽���-""x��v}"π�&
���i� 1R*���#5�x5�?t��b�p��<��MIh�t���n&%���Nh�kpp���k /XY 5䰘r��eβO��xps��l.{�^M��l�* a��� ����؆�`*	�6���]�����»)��I��hwe���0��a�N] ��`*�Enx~v�Rn��tq�kZܧO7q���Y}��9�B�- %����
'��"hց����kPA׬�9 ���{��GG%n箦�u�@�Ά���-���g@��K/gl�Cgl%FaW=�Re�\���q��[��)�|�Ғ7�Mn?Lk6[W]ҫb�iW��; �H$n����7����&=׹#������)���AR�J�RQ�d`UO��r��$�|v�V�o�l4a7܇YoL�i��첮��e�������t� (R������<����h�	���}��%�����N$B��'�ru��L~�q�~�W����^M�g-�H���p�32:
0����X��l;Ɏ��6��V�䝡��\����0�a���y���
*%�����J��I:�
듅 �T��`�ѳ~'Gǝi�GP��g=$�iDq��d>�����I@�w%��Ot��H�8r��<�ċ_e���p�g��̨�u��on�y�L�=mA{]���8�bG|e0o��b�[B�,_�O 1��6��i	uA==��溔):k� �AG_��w��v�e���fgcc�Й0R�Vӣ��#:8��Uez{ߡxЉW�á2�V�w��%ҢU���|ȡ`))z>]�p��G�g}��nb$�{��3�.,X�6:xN��$f�i�xe���]�n,����͖G��P�l��zuQ�:25�R��)�����Eg�����`����������X���ǽ4�^1�1d�z�L��,������+��f�#�0�2S`{jZZ����(�-���3�r<��_��"r�邱n�S�5E9�Őw��K�"I@.J� ��bj+Sp/��:04Tъ��ϰ�72*D���2kW�'�ګ4�zy���V/��ٹ�^ׯ� 409�軄���mO��E=G,.vC�j41K\�2b��+������>���T���P}���%Q,Y
b�R��Ԕ�����cPSȶdX��c�o�Ru3�b?άB��'UIߥ��p�w�˶F�}!�2^>\�Eh����Y9�<	 _������ͣc��BN/>��سW17�����srrv��pȘ�+���)&<z���c��6n����
�����QXA`@A`W	i�	EB�;T�:TXBPR�s�!D��a:��� ~�g�����}�=�\+��k�G@�Y���u��Nn9�]s�yGA�2�vonA���|��rF(���}�!��'l�rm�B&��+f�2 E�{q��&��ۋ~Mj�o˺?WX�@7��q3��V�� ����������Vj���@��
b�c��+<@-�m�Ėp�N4H�y*T�.d|6���
V:���nn+_H�\��q���\*;�E�C��w���?5c*���� ��ǧM+|@@ �/y-���M�Ha��"�;��	;�v��o� bf3�!�/�v
�liyB+�k�cU � %�4��q�S������5$$$;�#���k����?䈖|	��q��y���Þ T�7�	���r[��$lb�S6��5�.y�t��1���D �M����9tV��osW�w�.w.{=�(٢�_��@k�[�B���q*��x|tJMC���Bm���ZF�V��#�k	2�3����XĹ/He�t�(9C~Z��i>����� ���x����� �iB�e��$�����\�q���+��sN���{?�%+��)�_b�ٸkW���j:/�+(��!K�ń>�=��%6��0���a��&��~��Ϝڿ�� � ��۫����'��?� 1Z�*���I
?�؏��(ԭ�.�p	~~��z8���S�:�Uq]���^���G��+�S��ώ��&�WhY��=~��rs)�����u��hu�+�s-`'�.h"�%��W�T
��E�F�N��OGЉB��I��$e��П�$��dU��ma�%���@��͸�{M2��CPm�[M��){g�h�i��W��Q��@�:.qtT��TL���=vJ�_)�k.w/#d�s��Ma?	b�Y�dr`|�-��%q@�@9��kf�h����o�=�g:\�Z����Q����]ETW=ڔ����㺘%%��珃]o���|�<+/�����eQz��㛞~�ƃH�˵��<�Q	�ѷ�Ԟ9�-�U�='&��9� |�@՟ W����p�E�=�vhv�Tj,�ݏ�'dA���A_�S�c��Rt���g�UH�I��e�fݔ�h4�ȿ��@"
�B�+1��_�I],Fh�bq����
������zßI�HC�!��.ۋ�c��\��YH�ɵ�R� �#n������[���&C;�����mAپ#1��ֲ�k@fj+ЍѤ\�c3�V  Y�5��;���;� %�\~e�U�[�x��Y	(�����}y{�ѫ���n�[��9� R�l��FF�ம�a%F�z��3���sF�<׫,���
�(����+-��/Ҏ�|�/Kc_ov;��ڛpӧ��|`��h3E#^�ͤ��\��_��m��azt���.]2���t缴�mj��x^��QHL��(}q�UD��x�ɳe��(�yG�޾��N���_!���$0 nO~��ް.U���� m��/]��q���Ȭ����Xf�X�,�Zl�[		�\����>��S��Ijkkc����N%��������K{�(i�2_��x��ˮ���Ίt��u���|Hq,M�.Ӛ�9������� *xK䤜S�)Ub7V���a3�D�A��X����˨ͫ׷��ѝQ�ݓ���J@6�AOx&˿�#Mf�9!��yu��-��E󮯭�9��(����~	6\�k�'ٗ"� ���fs��V�8�t����l������<ɻ�CVj%SXQQQ3����|'�ml5<t�_��N|��YZO���������-��kЊtY��jeffR���\�J�h�W��̭K_`�\m���Ye�� �0 X���h��B�~�����\�r*�W�QW�܎'I����}��m���'�vdm�f(����J� lY ���j4�k���Bh��\�|>F�K���v�*��W�Dڗ`��5W�{�����ņ�"�����;{{qU�_����W��h��+3E���%tW�Tb1���k��#������_.���A~�����z}��io�y]N�OV2z+V�%�M�,�9�sM���A 
�� 	�~�֠8�6---N��Vkv�X�p	�s�K��U�$��⻯�6�.e N�����"%%-��.����T������\vz�!� h�Qh{��k�ϵ�˲y���� ��jۜ����u�������*�""����Ȏo^,8!��1r����5W��U�6 [Z��������Kz6QB6n+ ��#��ҫ6w(_��G���t5�7X-_��PWW7K�N;Z�&��>�>�\ᙙC�M��p��D�����-��i:�}�����k׮up_+2D�,?����c��D�hlUdd���Oz���*�@��U-�A}�SL�/$�멧�G�&���J9��ը�����mY��|e��쬠�b�< _�F����o�g����7���'�m���҅�O27�j�xԩ��>�U�X 6g��U���t=�-' P��ҫ:��.�~���U�΢,��������..���{��/���N�^�_@ @������<|iܘ�s����0�TĀ3̎��/�|�{-��w�Հ���XŚ��ug��nL0�j�/:���h|7"���ٝ�:θ������T؛.a7|��*�^jD��of"{�h��O����VV� �궯A��?������3Dw��(�R񸸸䥧��8��kP�?�7C=9����~
��: �u���|�-��}�A�e�!�<��0�� ����:Sⵉے�r�ܧ.����rv����{�����sN���[�l�G�tc��c����'��
Pe�jM<�ʣ��R�i��6]�}h�"m��T1
m�d�;�������L����}���tͫ)��.=�~2���) �k���Jn=�/(�K	-���o�Tf5��,�S&��a|~˻�B�7%C�4Í�P.5p��&$�g��UX}||��
�Dv.���C��===�8e�J)�P������f��Ѥ�b�ԍ
�q��_D��əW��m�����ӥ`������,3�'�Xb��9K\�I�����M=�A^����}�<�c��� �C�\zE�����Xj����=|����?K��
C�B�/��3Z����x�V� �%�����h�P5���ik�4+�2@@-��X��;!l�#���#?~���h�?`YF�����L��xN/Z.j�[�W��rF�ŭ�|nx�^R:m�,�U:s��̘�Xx=�����Gx�w�������u���bK=���/�m�T��8NC57����1>ᮁ��eu��\���>���>�ap�tw܁�,Tx|�\�¾}u��P��u444������`D[��;��t��C�;k��Ĭ�i.ĥ��-���@��l����g��Қv�#a�%~P��}%��>�NQ���o�'�O�p}mL�̶ۘ*r������u���PϬ��$��mƞ��� co__AnnЯp~(��{�6ŏ�Z܁�(e�$c��g���;p����b�0��@ 	խ�g]N%����i-[K��ד{ע��Mx��mu1��]���"+�"��O��:�<V��"�R%��yg�EJyUs���yd�t�ߜ��x�ĺ	q���kM�L4��[�STȳ{Z2����Rq�&+Az��������e�~.{��� �t?��ث������]o�
��,�Ғ�D�/@�b�W�ӟ��l��~E�C5[��c,�������F����ކ��������{�m��
x��M��e�k][�Y
L��rG�����w�~�1�X���8���<�~�XSǍQ4-�BlO���N�!H<�f7n2��X>1!�+����C��	�6���������* �%�iR� ���xyy��=(?j|���.�N9��g)��bn��?�A�dr�M|��n$�8� ¡��Zx�[Zק���]����C=�Xm@�L�
�g��t!�J��e�_���y���3I�� #,�
@@-3�����Q�ە9���bb���,�5�i���M28/���Tm�=通����&��<��pjq1��H�J��UXZʝ�����p���~s@3E:w���n\��C�߽3�Ϡ�D�vܾ�C�x���A!�ӆ��Dy��Z���l������l�ΝV��;`9Y{V�D��
�	�FZ��yb�h�{��4�(���M�~�����)@ 䓓��ի�� ��6M����	���O����j�?~|

���
 rc3��S r�B���1%h��{{�r��>���z����F2�w튑��@��$�|�q�������4&�SC�V��l�p<��ؾ��Rf|�Z���9�eu�b���d�~y���P��`�A3ʹч� �M+b ������D��y��U�ۏ���koEў��Be�y1�����=�Z���@���(�GXT�ֻ<_�K���$����S�
��b}����P������)���N�f{�s��
����6�-�V�	�{�`R�X�3���Կ*��s��i�'�r�T�a���W�u��j����s��RTVnn�H׸���s�j?����tܦˤ�'��9Щ3�.iz�ȓ���R��K��W�=���t�;r�A�΀�؜��5yd��w���9e�'�$��,�������r���ӭX'�T6����W�K�~�մ⹁)��m�MFG���"�{	�c��!��/�	����|�_�,lY�u�Pf�+j+E��ת�G؍il2YGCmB&6I��뉩1 ��f�bs�G2�	��Ƭ�E����TU<���^ ��kL[��w�CO�<	hȮ�r����p��@%��5$����Pg&�R�R��Ï�L5pGM�>X\Q�l��cW�k~���9�-Z.{xd�"�|��
L�`� JB�E755�ހ�nUp�s��D�L��I��zL�h�q�~ )���E�?@��	�
�ק�0���/0����Ⱦ��a���\S��Ʉщ��Z_�|�R��^�g+���a���o����mf���q\�Ts����������t|Fcͪ�55��FC���G�Xo��(yJ �1���IɃɳ��~'a���������	��p�M�r�` ��E�T%������,�gE'ם����
�@�p}ڴ����g��-��d:|m�'{	F⟧�jj��vZ���45}D���2y*��G*N��HFF�Y�%�d0҂���ϗ��m�lVE6�I��<���A���#����~LC��ag ?�mG3@̳����7cK����&�J�G!Ղ6�RdVJ�͟��-�7F�,��J���r��ϊ���������\���4��K���Ю>>���;+�V=)��B�bC$�0
�������)`�Y[���T�*b~;�;�ד*����o�#��A jU��˿�h��E`c�y��݃����\���rp(Yu��3�{�4�@� ���o�P߹S7��~?:��v98��"�������;	h��?�ʎ�؛= ɺ���i?���:�S�V�_�����b���\MP�X�ho���	��ӜS�� ����wG0r�sPx��~J�����+i�Ny�C������A�{��6���m�@WAe��So�n]#d�P�Kp�t6zx��>��R���J�y��H,�{Ǟ�d&�9�Q��hM|[�p�ЧBwsZha*�mmm����r���R#.v�sѧ��T�0�� ��ŮM�e��Z���]�J�~NuI��������&'��O�]#�b���eu�GZ���K/� ���f.��چ1�V�t��%�����#�q���>.����#i�V� R�K�~zP�t�Bsj���Qs�ՙ�D����gb�zz+-	q t8��<c������%당����_�jr7�O��
�ܘ��m6�t���0�"�� �g4�!DeƉo���u�������%��m�;�iil�>^`ޚ_��C�0IZ�u!��ֶ��6�뾚�.��U�k�BJq�	�,	�����>jض�F� �Mջ,�SMZ��K"ƃ?��U�"Ϊ���f=�Feo�]� o�T,ܱ����8�|�|�s�s �l�nE�;���=��-㍫P�����4}���V����!�N�ZG�CϪ�)��q�A=tWo����0)5F�j��^�k�/�N��A��6|y?�}��.���]3g+��I!��G� ���d߄��& 2�d�/���}���3<5�Nq�=Q%Xw7�8�ٛ�w�և���O��6�
��04���oBB��	hiE:��_Q��ʑ�W�Dj&=�W�%���q�2���ߡD�9G!9�2B7�D1#EW(���~�� #2T�o�	܅�
���M9��!򖆏���I@^�S�ݏJ�Ee��M2��7DT��A3���հ���P�/q �`�����to�\7���:r�aKDUom-�tM��rk�̖��:L%����
 ���'��'rF��/���u��Gwɤ�]7l���zyii��A:& �ol|\^ ���}[������/��PNz�'�<@	�p��/���]�:C	p �c��GCn6����~�v���xI//��|e9`��A�P�j�q�Q�R� �����%6�s��gz���\>�txP>'��	D�4yy���cW`*���ꛞ�w.�oI��TP�=���h��Z�D�tYHA �J���*_��Y����#j��'M�->c����m���V�����G��H��Zh5ED
z��м��˽����e�e��ֻ�%�$�2����2W��&3J�CɇP�E2Z�,��TBR��uIWO��S<�������ff���wP+���ܷ��&�����s�,�����2y��w-�x���W� �]�q߆���jƋ�5y#;����o��X�_&$$,����0��o��jV�ag��@��5�[�
��><q�D6"5�$S[ .�ᭂz&�T��o'l3~���$���R.�����XĽ	�T(S�?�j���'��!"��>����~���:9�'��о�u~�*��[������]k0➜��{B���
9J�"ǫ�����Z�����.�w��+j?0�ΰ��o�@P��|VΠ)��p�ky���r��wtxSխWW��]���X���r�mm	@�QA)��Gc�J�#W{���~ǸC��&��'n�8�����U�8����-�"r-�{��׾��&��៖�gҬ���r�nvY�����';h�=�GYZ��Ą5�D��$ "	Ll�J�����E�
b\^�:�n:������Q��笢���=��N�i��33��z�>�ی,����,)w���2Be���;�_���@�^s]���dӿ��W�t	or�%��C=�(���q[��蟩p�o�C�lBb���Xf�%(*(@�����m)	h2� Iy������l+�"�گj.O���ꏡ��S��/<�S^ {�l�U�p��i9�^;a�#����I�����*���F	 -��1���;y�c�Q- zɧU2|�5�1����� X�&%%]��G�-{������m4]!����R2<�_���dQ/-�$	����+ ����:89�ػ��� ���ɛUu��h���2ޛ)x�7��4v�C��������!�?ۡ��3��v+���\wu@��N7"V�|��Q(�u\OR�t�IB��Yf��0�"��?��$P `�Ag�7Jo����I(���B��V/�	%����>R����E�6Q?#n��T)�o����|��1Ҷ(��6���*�sobW	�c�*�^�ܣ�3���e�<'p���aM?����bW^l���#���3�S�7�{M�ԏ��݉~{U�Pϕ�V��n�0G�ޞ��C০�{����:���5�`�K�Fj�>�])�n5��p8��/������%6�* -w֣���,DS�x�+.�G��E�w M�W��e�MJ��Q���.�(�E��w��ם��!�����-�����	hy���l�;n'�_`nN��ןN�6(���GD�<�K("j�_ ����W�;�ƅ���7�|u��u�5W*d�VπTw-1&S�p5�P���ӣ�Z%0�>e֓�?���ho]�+ ���/��AOJJJd� v�8�D�JN+��[Xu����9[U7'�g�.��&܀'�h(��_��|r�б8m'p�T��=s��,=/�M�<>@m,i9e-�l�F��ĥj�`���Z�;�]���dVc�L	��W���H���C�\��˳�#'��s��y=�+zQ�zg��\�/	�f�s!�}8�o���Z�Ǧ��<]�u7S�s_��'���O.���եde̬sv��eX?��/OZ[閨�ϴUWd��8SD����(�Y9W�ڡ�h�����
�8�\s��Qy�����dd^^�pZX�hyOr2m�.n��}�Qv{�Y�X�ʆ	��o���h�r��:����_%hԕ*On:�X��I��^���+B���8�Z߂��ƴ�J΂�u&aq��s�!��z�(���^���4����\:P�R���W>��y�/��6j�ebbR>�f��Ps~�Tj9�~5��(:�N�����ӡ菟b?~�Z޼��D�Ip��bi�N�"$��߼�l�s[h����>������TP���[�b�4]���X̄�ƠG��vla_զ��y߇�'4.E���?���m��.��ژ����*�z�N�(�����c&Q�l��9�:Z��&KT~T��1�u�f��|c���P
�-�������+�=vJ��c,���dTT���	<�cy�W�R^���yj�0^b&¥3դ���\��p�YpEPh�q�6�NQz���*���&�#>11{xV�CQQ�������On��#,L��������"���´���|[r)���������=Wk��s�|�䭭�X��Ӡ��96ぶ�4���~���s����)���1t����Q�t袰�>>��呷�/�/{>�B���s\8��gs؏gR�3m7,�)�F�\��?���i=�5X� �3� ���Ne:
�/�m�Th�4���fN�	����E �/h�nz�{^�7��߿_?�!<����ޥ<j�}����NY�'C��������<Z7��>A��yz+D]����9
������";B�~M�Q>�G-�5��R"��W��7AǦ!����<��}�,��g|��'|�V3���o�i��n_o$~��5��"����ji�ٸI7g���_� W3�`~ۙ��?��B/���Y ��a|�XW�݊T�3��<C@�R�s+mGyD�V+���s��;'#�����{��/����˨F�\RRצv��h�Ǿf�--,�`n�`fR3>�2����A�+47*���՗��Y�L���j�N�,���{A\/������b��}��Z
�&�u�� �ֵ�����1G*)+#���L��X����}<�Urn�͈p�pu,�sy�VXdW�L�p���&�����t/Ĉ<��!�W�41��h�z�tX����	i'i&R��Y����h�>O$n��)ؕ��[3�jg!*��د�/�@�w�G���7�.8���	'U��ї�46��7K~�[��.����ؐeP�f���	����(U׬;����潴����}����4�'<%ic����/R|��K�[�/��2�4�%������t�?�-���֠v��2��ٵ��Ղ�C�yg����Y6l�#خP>��yT���V4�k�y�4g&$5G1��ѷ����d�E��a:� ��?�Xo.�8���9�M�z�D���e��NP�Q���W(�0'>.��į�SJ揮/=91�/tO�E���#GU�J'� zk�A�}�߸|?jz�����z�1GFFf`ż�{��i\��R��Pl:=@D�����k���/�~5u�N����V�T�;���4�=�/?�3>�.Xj4~�ߌ�"�L����	#v�a,zsb}���9���Q�e�JE-���1����u�|_��3�֠����������	�6�$�?I���]��+���|��u{8�����K�T_�(�fM��ҋ2'�d-l*����Χ��WJ���ti���1�<����(jV[G7��m�t����o�(�<��9ڵ�nh�ʏNAn=��ޕA^�Dlu��"�i��F��j�~�3��|ւhKu���(Y	:os�3�5���\؂�$mr~��I��u~N)�ҳ�I=�Z�O�7�R��I)��/���b	�+�M�����xѫ�X�,?����ou���LB��Y ��ݳ<f�8y����L�*�	a�fqY��fh��kUII�'Cǃos���?X��{�"r���\�e��	�sݴ�ŏ[�d2,R<�O�MҒ�������t2F%{'�����Y5Y^\|p��7u�3�鿯rw�� �)�����.�?���,�����DD_�����CR��E��b�w��ق�eZ����Q�Yff&tpxtT�q#�Y�
�M�����s���<�{]�)H�hyK�[=���6�]����y�lyg>��:�|-.<C�%,����t����^��E�I�R���49�,�xd�bO_Bo�e�@Y�@�;J���}^��@�J�i1��^_,F�i���Z�i_c`�Q�`��i�(��參@\k���QZ֩���Li��]�{dx���<ϔ?�%�ޘ�������9�Gd��	b�e�A�s�{���(�NN��{y�(�a~nnGu�g�J�P�����[�)�߆��U����3/MӒ����C�yQ���)0���I�b\˶�*:����KxXB�a%�BJ��NS��V��} �R��j78�(4��`Ek�0���Q��l���{E,�Xv�v�9����[	����u����:~����-�e��V� �5�9G!��:�R�o��l�_OT�:��+����Է?a0�
��b�`���
a�������:�b`Cd�A�L'LQ�E��	9���+Dr��=��[&Vv(i�2�a��rL��6�I�v�}*����V�s���h�S�W��q.�	9
�!�iH�u�wƵ@S6���G"C��#H'�G�U�9\�Z*D�`�:ۯ�z �M��ٝ{�K��RXZ��UzkQt���X�����,�|���K�[��N���cKt���Y��
L��R��A�uO{�k�ʁ����d:O
�9^g��6����0~�}�I��$�����Q��5OvBGQ(I��""'7W�\vF.����xſ��ۡ���&�`��~���~K����?��3�IN^,u�Dz,0��2(�ĩ.if�=��e��F�?.���J:���o��BTkP��}#�lOLa�w�����p�<�	��31''���gW�>��9�4l�6W�PX��_�et�)T]�?.%'P~z�cdd$ݾw��y�s�+��n��6�����Q�9hP3���� �����J��D{ �s�;�A�K���Ax�Ό����{Ή����Z4NCV_귨�%����	���xG[FC�-�����6������"� ��	&�������������U��!��qv~��b�#z�l�����p�n�,;�߹ j40���c�70X}�E��T��vy��+q�t|0��L |�W�/t�� �ݴ�D�20���t��þþ��F������0�#�r��;��F�&��'�����^�]�a��U�H cGb�_�R��]5u��w����#�宓��f�C�|���/��s;�;#���L/?��G������`�/	��8�x�V��%� ���mv~x=�C�$��4bh�b$~�ޜ&Ee��`*���9�B�:�9�^{ˋ��e��V	��&�\(��k�"u'���u~F����꿚/��Ө4w��]�rV����JB��j]F!�����;VW�T݁Հ��!#d���?�����ӢGK�x��l�x�FX�<��i�3�#�yx2pZ�y���P�*p>�w�N5�z>�%CM��GGu���Z���
ݍ}y*��i&*Fw2(�[ֵ95翉{4��\w�w�牊3��z*��ӄ��۔!�$���fuN����ca����lJ����C��+������C�"č*}�Ӏ����������uq��)m�a��/�jg���j]� _����dq;��B�D����J�ˑ�]K�]� ��Bi�D�.�;�����vK��7���>=§��Qc�^�i( 3���5>��1!��m���׏��KU^)B�y�
A�\���.�Q�+���F˳������,Ӏ�`��ո�/_�Q
�J�~�\����Q��]|<`ݯ�a6���3��G��~�$ϔ'_���u	:)�^�Y��x��We<뮾��jE{��>�.���K���5R�Ni�����d/uz�7�=M�'0j6��oE��փ�f�r�؟?K!��`�~�m	OB�N6��/����=���Lu	&�Sz��w	�M�Y+sQ���Q7�b���)��x�$%��<���V\r��po`غ\]���bk�ͱ�Զv6�{�X�ɹF��k��4��t!#�tlw{�enș'/M��JH&@��%o�|�9�1�
�Ha�m򡦦.X�[��8Cgĸ��;�G����4ΘMIB�+��jօ�������te�"�� �ʔj����s e��5C���~�����9h5�x�M�F���>!7T�^��/&�N�e��$�|�q+,��?p8<�__��p�/4Iȁ�82e" �c_����@Y��t@p�$ә2�, ���N�J��YXU�|�4|���B��BÑ�����PV��tr�����,�
�9Q�lY�õ	�6��)���B'f�$�_Pa�4����f��ù�oX�h��[��v��]B�JP� ��"�*CθX}�ꃗ��o��w���٨�^g��B"�6T�;��t>5_���r	 wyΘǿ��%&"0�@�c
k���쫸\~	�<�0���a�'���3����_i�N���o��g�X4(��+�!�YM8���`ζZ?��'YEst���ѕ���9���+�ش��P!���6���EF���H���~M��*�p8tt|��@��^�wh"���tJop�*YN)���4oF��ΰM-���O3�`kF}9B-L:���'BX�5�S2i���}�\L�ŵ���6�2Gկ��}�J��^p�P�A��Q��`�{���*W�v	|��F$v���Ȧ��^���f_��VBk�T-��h�Vq[�0������ ����[z#c@�G�ǽ���d<Vˏ���۷���]G�0�D��*ӎ�/O����:�=sa����%u��(����~:���p�x�
���**�!�
�m��d[��[����'@x�>vW!"���
_�GF;�њ�6��>;w��kw6BP����M^��bXM�p���f��I{8K�KƹW�	9��GvP"`W5��p�p��y�M���+\@=�>a�6����.}�eX���%ӭ���Ac-����/�qo}[�̸�&\zV�Re���f%�k@����^p����E�7��2�M�}�)/B������w��{�>�ӓTh�=�mR��nge&������o������!@��pu'�|�-�w�r"�,6�
���^��{��	{ƨ�/�?[W�*W�*��(�P�:d��?!�� U�p�?��3?*A#$������������5���㓅Z�����]�=l4~�ݔ�/���⮮���ץ��SL��Д����	��<\���%���4Ȩ��`�/v�U��\����~�0���������S���4���W g���eW���G�W���+7ズn.������<�į��-*��rg<_:�:;�L@�����9�`������U:�u�L~�u*N���������x�Q�ή��#^��u}}QΜ�+|��z M�u]w)����9^�� �hɂF
u�G�|||��YlH��P��&֚qßU�UW$���u�=�3�1��h�R����@\{��gʾv��.���D��V���B��W�Q�S]@򟟐�J�G�<��&���6��Fю6 sU� ͣ<�3a�a+ U�E�̴^%%'G��w�h�Y�R�&&&���P� ˂�&���L�uN%�ӳa	��=�=l"^[2�ΣD,ഏ�Kh0��z*.#������DН���8D�Vsue�b���meC<zn��������B }?74�7Л�J}L���1B��H��8tw��o`�V@�����WBэ֛P���v�\�84���#ګ,��*���8R�O�9�{�;P��{��Sl��q���v×�5e#_�(/,"ҭ�fn.��>~� "=�(���X�:5�����4 �)Ӵ�����H��w��nŋ���dʙ��}�E��Jko��Zr	��$ ��Bm�����e��NC.���v��I���ț������W2|��n�,��������%�UPm�< ��K���r�j���[�Yʏ ] �vwיv��,���I���I�i�O�|�j<��^1�Ku�A��.s7�̌�q��$&nT��8R��b9 �	�:;%�vQ��i�o�T#�9
Z!Ǵ�ܲ>��%έ�o<;�����f�8iy�W���ᖂ���T�T�f��+Q�U*�����t�:@�#���W!�Ζ���X;��-����:��hHd���k�3��S��N�ﴂ��*�ȿl
�Z�r�G;����q3��������������o��v>Eu�x7ǚe��}m)��E3�9Ң��ͯ�Q������ps��?6�>PfVJ�������X3nO*а�r�CM�5�zB$,tsk&��'��8����G8���*uh�_ٺ�&����}�6m|�Y߃*tQ�{�Nrv�"�3�!%#���)�I����6�.�,Q�&^�-������̙��Xe���lk��==k	))#����K���m�SD�q���՞omgg�k�No�:�@�˂%e}��->|	��i_Ӎ�С��6��H��о�|$�8M\MA[����x��G��@��E}T�-�Nq �w�3F���<K������)1^��A5='~dA���2o��&��ع$is��<|F$911a��k�B��c�T����!�JHDD��0����d�z�/>��%���$F�k؀�� �+?x�m��ۂ�x}��{�tW���j�C�Ru��/��?�!������x�B@� �����mZF��j�&���S5j�X"����Hڻ�^6Ϻ�������$g����at�i��}�UTF�(� �@��`��]�q;U����B��{�����i����ǖ���{�Q_̣x�߬��>e�*'���΁�ׯ�?���fK�ק�
���GE[f����$������J@'#t��OKLhDj�Ԙ��XxS�ax'R����Bw ��w5hF��=&��ݬ !	��5er�	�H���>�H�2��\�\��	,Oη�9ǁ�+��~�8�DT�T����]N��p�+d-z���P��)�;�GNNN>�4�];�c7��O�������6B�B�|���Ϝ?�bl��L���g֏��R���^9M��Q��I�uKV�o�+	�2����u�����E�U�udј\yg=�Z�k�l���pS����[�l��,��i���_�������Ϙ	Q��
�����<��|�4�S�׏.q/.-��a�I��5�R^�09�	

rX����mf��=����-6.~��:[�GM��n�.dV:���談6^(_�A�7w؛��7��%��V~�P�э|��a\2��M�M�v-�WՖS;{�GM�-	U��0�Ǐ�S��n޼	��kr��>���ܕ�o�����|��nC����q^-�x��?�F B�-��ݰ�.�,dH�+J!-#C�r0鵞o�)R.ho��1��(Ǚ�D��	q���s7/�=X�pf���Y�CE��g_�n������j"w	f�-��|r���,�}wL��O�6.Tn"�|�J��ի��_��Lk/
nŽ�����ucœ���xz� ��tu ��|{5��],���[�SL�Q�,��R��*�z�m���w�E����m
9������O�H@5���� ��&
�K��eX9_� �-
$t�I����]Y��5�MP�
�E=��{�n�8��Y�C�^���ww�e4��bz�'��%�+�`ħv<)���eW����=�g��ym�>)��$����faa�{����Z{���p����.���/vTX�* �m�����ָ�\�M��>'�eJz::y��@�Px���/.��$�>���t1%��k�9X�J�H�Z?�+��^9�{� Z.F�J1^юS�V�������?br��3���b����ZՇX]�GF�BG�᫈Ɗ�e�v=����9S^U��G	�D����1������f$.�L�G��,]LO__n�]&����\,\p0[KYc�����;�k�a�U��egg2[)����w4BK[Z��x�:�\�ة�_9�V&�Wz�� �?e#�ۼ�W�}���dffV�Y�A���1�$�eg ����s������;䷉�)�2>�O������L	)�We��ލ_�~o}z9K*5�2����>%f{���Û�C��C�:�89t�99i�x�j|Β+��
 &��^��s|T�7�sX��ܷtt�䫕,W�,����) l�t�X&S��:f�������>����{3v�5�:* �l; �y�) S�����$ԃ���2�����u����T�j\Y�r>�n8���N`��Gj�K��v����~#?~|R˿u⬣ma�p���8��!�4F' �n��}�T�1.�L+��o�aWLED����Ǯځ�		I�zh������+b��{/b'ȚڟK+�:\�Pܐ߃�B�c\��K�Q0�~�(��a�5f[�IG��2"��knm4�l�K�5&�b_kO���j�ʁGӊzj\@\b�������8B-�����~0����sg�pZ��_߰���IM�
�m��v���"\d��!��2�*Bv����lb'��4���0�[�z�/m���]�q��|S ����MB<�m���+<�w�������ٶ�`��n u��l��ӿ ��!7��q#`�ç-��w��;�g�G'��B�V>ՠ
ɯ]����rB�33�Q�!�]��7���-�{{	).�^ϙ��{�o�q <� �İiC��|��<h�~q��)��]��lx�?���Y��2sD��A�e�Zy4Q��@D�R:���d�z-r��|��̎ҟ:U�(�}��<�>vs3M�p�#/��sKˎ]=�b�2�a�����V������gcu��zU�fvĝ�!��� ��k��Ŝ	���_2�X��[oF�4��e���W�{�5��ƨ�?2���7��dY��K�\�U�?	��WW+�=ob�4�M�� ���N�i�e�g�#��z�U�D�%�2dXO��l4�pl7qSP��j����֭�o�p�R���zR6f_l �ӫ����� ���pO��]�T��8��#�"��j�q�'G�f��+8�u�ʘ�ړF��0aaaK^�J�d��TSid�p���޾���SzZ�M�$�j8����Hz�b�+Ā�x����k�����hxbb��.j5��Ғ�SU�UĿ��`X5��oߤjL �U�}����N�$d��u�aMfM;ꂫ���"��T�w\Q@zG�J/�C��"������^B���C@D�I	�tBB����~�%?�}w�9���}�s��H�UKo&�e�Ϟl�}���l& $T����e�TY��������9�Qd�̯�GTp����(C�\:���Qz�q��\�cy���ّ;����ؼ�����%��	:,|��'��CoK�)��pD�j|�#J���jq�:���[gQ�_\RRQ\www�&����2~E��^]`��!i�����2Gޓ�f���$�g啕�_�̅�ea�����a���_ �XI��]�u.�^V��[�o�QÄn"�I�}��N�1�� 7�Ã��l����nTʲ1�%�j���Y$0z��_#\�cC#��H���eM(M�0����zJX5�w��s�'L��ҏ����4�D0���p�Q��@l'	H���R�ԢJ��o��q�0*+ݒ2�!i�$ͼ���t���/D �Rew�.�+�>(�����'��t?;���\�����E��z��bf�߹�08j3v����� �CxWb\gIH%�{y��N�XD�o_�~�<}�9�{������kc�9p ��N�$�J�sC �4;;`��,��q&{����z�<]䔑����;�����t�E�Y���P�SE��ڽ�ܞƋ���,��O��ݝj%�j��:C 5��p���7�VҠ�L�a�&&S����j�T'n͜{�\�����hZHXg~f��hg{{�����I�f۠^��h�-��`I�LC�s�� n-d߄��T���]pdI�|\��N�&/`���_~<���~o[��ۊ
>|�sV�E�w�τ�uL�?}M�Do��:���D�9�������ꇠ���I�����|
�K`2{��N!�@����;�T:��..�����Md��y"�G>跷�2�ʋ�+볲��%j����c(�1W9���>���������p�����vN��Q�h�����67���0���Oa|#Y߆XܥV�3�4wE?��;�QMoo��^G�pIn�_�*X��;T� ��A7����
� �C��"���3g/.�d�Ũ�� �87��ep�b�&���r�^����/kNtWF������rkRcufZ��c}���[�+�g;⅄�r �Vxs�Hw��P�\7q�o#�jܳ3�V4�F��6sA)��bêvA�*�b#�&V�����e�D�4�"}Sά�_4:F۴s�j�d[ĝ/������>4My}wf���9��4��Ѩ�����c߾D}����xM����Pa��-at@�gyJ�\8G߂��1�o:�v������u��|��/Guս�S�$�aĒ���b��B�ޞ�~�p��p�J���;]]]�׽K�|fq�~�b�Ĭ�D�N=y�~R@��{
�H)%%��� �wG ky�HɌ�õg+9�"?߮�ʂ�˘:DY��#�a*O�Id|v�Ī�q>r�U^�Y}zNEU� /O��<Z����k��p�L*_܇�![�����i�I 	�a�gΎ��4�0 A֛�Q�WI�-qƾ�&��w!�8����5~D�4�*[�NS�)r����z�Ɗm��g�aLӑ4\��;���N+s�� f&&'������G�^jz�.+����mY.dGgu���!��Ë��o@�r���Yn�^�}��_�v��U��$K:C<��nZ7�ҴP�g����\�Ipț����-$h������� ZS�W��oit6�9��4���;X�N��ϷsrR�R�])���\M��a,��c�eQ��9pt��p�k&%w��yڽ��謫���ۜ	5eX�߄cll�r���AqBJ� ԥ$��*D#��?�u	@�(c�I�J��e�����S��q�5�{B	-EA���'��G�l�O�=mH��U��G�K>���a��@`u~�n����\-�k{�o[�4;��fu=?k����l'|7T���Π�����Tϟ�f7���2n��˵0kkP�'��2���&�`��uP|�Sv�a�`��]�3u,�ք�@��\�� ��2t�w-l�lncn���d��4?p�Ls�C��s�!YK�ok�WC~���Csq���g������`f�郌4ws��EX'»L��ߒV�n�C�)XE(�)����e��nU<����n���ɯ�$�-���UiUQ&h@�o<�B�eEmzU��JRB���`	7�N�_;Xa��8˲�#�1X�]��LP��z�/���e�r�I:��Xݗ�qPe(+y5j��-q��]���Ď�Y�d�G���
��56M��}�g�pU��B1t��&M���O��t��e��/0X��\�:�!�"&,-(�8g�j�V '?�u;�����+�1�݁������i(��w��V���u�G�,�+�#������Α��ϑtk���j�)))��46F�cu�ɇ^��݅��1_=�������5_)��p�]���7`���V.���dv�޷�P�(]�}J���IIZ����i6a��. �����*�������a �����������%��ס|,��ϖ�ĄI��������e�>��	�i����ЪR���4|�h��
�ņ�}/�z��@�P���4����!�Xd1`Кyʩ���pY,!h$�����A�w��Vby'�U����g�{L.y�����H"4�%�����ydVV�����-�<��:C(bG,�ߣt��4$R�jj��C�(��Ih*�Χ�����\��bKb;��B\o����q����8�$�p�Mi�Aԋ�Bac=Ϋ9}6�m�7���["��2c�.\\\#�pC"E�6�=)���~����+p��kY�����<��@V���["�uj���R�V̉�x���+.4�vd�-���5��L=n^"B����GFB�� ڌ��54�T����<"�`����⧅z����?��W�SN�<i����Q�xr�D���>E�Gj:��Q��l��ɭ~-�rhI��L����N;�A�ѳ��8}������h�{u�gaN���A`ͳ�J��ޗ�TƵh��i��X�(�#�s�E�-CwP_u\�1�YTz�Mq<����/��n���>A��p̈́�;�++g;�(w��Gி��ϧ}����Bj�Wb�3w�}Ԡ�Y6!����mK��
���1�(:�3��J�b���t��b���3��XIUG�������~lnV���`�wQ�B�if]�h�~/���D�i̴��f��>�Ӌ�`˄
�|Sw2V�����x�Ӗ�F	]}iV�ۿ�X]xS�g/�<˚��nM�
3Bl�`�w	����
5Y}�h�sX��8@��P=��׍�v@ެ	�8,i߾�H�=^s;%����k
�}�Tu!\jw��%���0��u�]g�d���	`9W�w5�NzgQE���Ź�$C���N7��rz�BmH��q'zdS[��i�
����q''i�G9�����<��ı�\.eN�r��X�W�V�.i|Em�#���c�ӵ9��^��)�)��[��V�� �rP*�Ø� _����"��^���lo8(���K�����6�f������/�2|���D~��>�Xw�/�8üߟe�p���=�*�%(-�����궐 �V�,��bF��`�GDK�ߧ�jN�����>��l���åB���1�u���6�6!/ �_�gB	�\�3����źBbbP.?`ٌ Tmh�d�"z�F�3����ln�i����o2��'l����߯=&�ӧ������2(��.
}%L�<��u�a7�n���y��ꆧ$b#X�
�ߚ����<���([�<�+�s�������s��_�h�Tt�D�K����*���*���@�	�6���R���k��O�D����C���J��l��:<\�\e3ۑe�AX��Zf
��93sss�q0N����"�	Y�U����7��i�W)�������0Tj�D  py~�#����G<�ħ��e7�m��{k-�|2l�,�`�Y۴�zTqLk�p�G(�$���4n��3(w�E�5�}��ٚ���q	����MC�0F��Z�ow��A�۴@3��QZ��	d�=�FE]z���v�=w�� �رmB�Y9y���P=_&�j�P�������*s��W%S��R���uwG[�}5J���� �ѣ4� ��v8��� ɺ����\d����Uw����GeJ� �(h����TNS��R��%��Z����A14<�J�ރ�K�>��vZ7�S�}im�g���o�ӣoxE�z(/Dz��#���ɸ�������Z�J���?v"j��(��,�*�<�τ�R�7I�v�1�>:BͩJy�m�.�vԿp��[%���AC�Ž�4=@��_w���X��W�$��ckҀg��c����ts�?�RT�q�lT~?��p*=���w	�x��R�s������e�U'�@�]ϴ��$�"��[#���w^��<�ӀQ*��bXz}��ߍR�⢢��W�N�Q+�b���q`8�}�p.����[" �(��f4L}��\�]��U���M"8 �w��m�֥�:^��k�F7�)�+m�ėo���Ti7K�*2A������~�#9996$�ٿ~��'�P[�s+��;1OS��ۃ[S���f�R���(�����| a���]p0��^�Sк��!���4�cM�Z��Kn����F�x�+�a_��IM������\�?#c��#++�_f�vE�����:���x��ZE��.��J�b��DSW	@영��w�Y�S�u��Dg��r2m��au��������Ss�l����͜��,�М|?��QSV��	G�e��[.��J�+ԓ����A��}1�Y25\�+VxS�07���a)\d\���Y"��.g,T�ݔ ͍�YY\D֙���ct����v��^��x
�,�#���xϱs�OO@����ۖ[��{�5�-;G�����E�i��G�#[�  ���y+�Ń[h ����6glE����z,��N�_%��������퇁>u���-z/3��sgEչ-FC|�eУ�U�顱��@KA��g{ٹHs�t���Q8��61t�6ko$�rZ�3� j\�g�V�Xa�$��@����w��t�w�UǊ�����Tˍ*� D ��}s�]w��r�G�F��Y$�*����0#w4XL���D��.�X_��3�j.��d�lE�{����f�O��hll����-pf�:��H.�fl5��8U�����,sG?N۠fɃ
�(�����ClGױ$�^x���؏-���;���f?��g-�OKJ�r���nm��H���i�[ڜ�vV��ꜱ�2B��F}0޾)����ǁ>I����|��r��ˋ��%N�ܥ��|����VP��1Jl���V2�-� #޵,M��օsk��$��1�)��r*],!������	ɳ��Ϝ9s�2hVF�D�ߑ~Pp��Xe�i��]�ez� ͓�^���xs���� ���pW󕖖�D�KNA�;������g¶���%^�&�?��M������w7E���\��  +ц>*b,"�#��\��Ãj�3�Y��c[.�b�b��?��������v�wĪJ�&K�j��F�'�$��TJf�6���c=��&�kO�.������#�<�Ӛ��������+��n�����.'��O\�������muDĈ���!�5�R q�D"�
}�[�`�~F:Hm��Q��T󶠧�Q�,����WF��c*J\�ۈRk�b��z� #�5��YjM�̃�ڞ������4����I�X7ť�$[l[qҞ����cb�*V��\UĔ/��u���RQ�'�eE�}�����˥�q�Ôp�l���&��G�V�ǲ�v��_|�˭��>5����ig�i��r���@A��6��	*N�k�+O��t��%5k�Pv:���"17..�m��H>��-,���M������9�?��/�병:���e�,�Q	]�I��k'*�,������"�1��/K��	+xLɄ�� �7����m�W��8���^�mm|���������x��P��q��� ]��|iU.���?3����=QNb��&U��H���6�J�Ӂ�3F���xxx;E&��bw�:o�#I��'�o/|�0}�/����NC`��nٛ�D����\�LǸ����'
�1[obTbq�;�{[���΍b����x!\ _�hl�tE�h��:��ٌ�<��P����7�gM�@�2�S�p�Umŉ�]$"�^��ޜ�����l@&+**�	vn�����饥�h6s��~}���?z"�b�4��2{12�7/�|������E�3�=ҳ���B��a�i���w,�(-��7�/����L�`�kz�{x��##KvZ���da鋬<<t�>���ަן��h�.-@�:�~*�ʺ�o}�D����*�rz�k�}{�y��S�*b�"��HU��I��W���I�*��K�p�ƀ	���n���_hg J�仨I�}*�#�����4ռض�m���⼴����
��ws�r��5��d2�� �۬�?�c�ҕ.��L�X�)I��&�:>^��&��}+j�vd�L����Alŭܖc=NWFO�#;��	 r�q+k�0�^E���2��G��񟐜�����X���l�;��κ�4������W�|��'����lB�#���.��1-wH�Mէo�˄<Ѐ�N��!`�W��NU�m���%�F/[&�BA���m��Qk Y�>�彄���HV���k��(+`��-��3"�������`K]P$��Ь����D�ؑ��10���iZ��j�">@L�&�J.�����C#��{����;��ڼ|�yP*���{����"�	��%�Xׇ�!�e��)���k����*���أm�~��������V��D��Ϭ�N5C��wv��3L1K�_��x�{UW��S�ȸg ������5�?��ɘ����#��\�z��-�I����=�@jA�����É%;L�������)UI1|K�����}�9C`�~&%(�0�.�
�ٚd�ܚ�)Y
T��~��0�"^a�>�XŜ��@�%�>Q"�J�B��DL��ԙF����|$���P�Z@���76������)��N��&��	n�Q~*��￙�j�����|�)�Չ^i����:3YenJ��twFv��8C������r�`���`#A�u��#��/��J6��A==!A�l�Cx-���\�i�[0� ֥�hv�j�'��x��ㅟj�>�9�rb#�&'���Kd���K�=��O%[�A�Е6�5V�͡&��Z4$�i�ո�l�ގ�+W��-\sDq�}�u�p�0��V	�co�Yvs��m��5�%ٸ���I��0r�D�?�����b�9���Y�� ��bccC�u�w�˷�������TF2��1m����B����ݐ��{4�ׅ��">�H��p��N{{{붡ܯa"�L%⬼��k�J,����~�1$����^Q���WӏQ?Oq��n1��'IڷI��o��v{ۧ>�h����鵒ޠ'��E+A�#}$���o�����߈����:}pC�}ˉKVە��9-�裴9�'}�1	>?l��V��H�YHٰ��1�S@`fo�}�pQ\|<�䀔�hl�TxE��;}x(;�B�O$��L�%�?6�P__Lʓvbz~���H��	��0�%�j�.���`��7��G���1�|�����"��$���)����1�b��������9�s	�o
�
��k��?�Eyy�!��J�|���ٟEl�r^����x�sd,�n�(ieeu��;s��yI�T�⦪��>�۾5q����j�$����_)�R��bMդ�>�\��;��9^N�Dz�2;�[�:~:��}�����&  ��|6j��{�5|��>�dlYq�4���_%�Oݕ�Bg�o��́�S`�<K�D�m̻O}����jxX_�36�.��o��q>1)�=yO�S{��4��I��SZ�*��)@)wJ�rfOn]�;�g������)ԁ�q<���@K�$~�O���?M���|D�0R>�!?5	��Q�%j����Zg��{��<�\�[P#jq�-amN���U���56�?%F5/}�( l�я=����D��	���`o{n_��0J�s�|熹�IZZZ��,J1'3�b"�������� Q��r��g�K�Q�~�RLO�TW��)K�z��&\��@o\����U9�|6�+�V����ݲ��d` ̊�(< w�D�W��t�G��]Z#
#���ЃT�w��_i����Q��Lz~<���J�=ҵP��'�����/_H� �]�7Tj���2V�S��L���s��a|Y�ֳ���VhL�uZ�B}���s����&{�#�^��D��`�5E��\����Tsyx�M�.I�|1�s��G�*R�ȸ�bWlm��������&�j�z���44\ש
�q���,@����ј���VsW3��V�ޭ&W/�X?5��0���,%&��(���w�h���)�M}S��|���;0�C룚��p���ٰ�����{����K�+�z6.g_	�HJ�N��)sL�0��~�8������=�O��i�,�?���988趷n���AxD���|����j�������ǎsչ�|�)$��B}{Y�dK����6'|�a��(��b���	j'�a�;U���ջL'z��M�yRP�+�l��Q���$�S��lu�vP��r?�G��#v(�},ܡ5�9��O�U��MA�
#Jg�b7��Q~I�`���IHe�TS^>�Į.����ܽ�c8����nc�@<��L��ڇ])�Yx֟ߴ��V�W�\s�+J�:b��vq`�d-���
�_{��rt,pK��jqq147Rq3k�ZS��$cAN|#���~�|C���#f��n��/����SE������VHI����/�2X�菝%{t�Z��L�1c���4�_��vF��i\�s�����E��Y�͐����
���\xډh/�$K�U���iERu���S�9�o�J����vNjy}Е���\��ܐ�"h��$�yuQ&����6�1w�j|���>�i���2L��7t����^2��5X��i�k���<]��E<��$^�,���Dj��o�d��?�Xt�����%������[�$�t�X^^�]�����:�{P���(�N��>��#j#��I����V��G�½��e�Bd3 N�=΋8�p�j��z��Q��iaa�;�ș�L��}?���4��T֯s��t'�A.�k��������҇��p�=D&'2�����Ya(��S��b=������F�7���o�KF�M {{^�	��)����y�t��g���{Wk�>.��@,<�l��Z �4��f�*X�&�P�9������4�C��z��\}�wNT�S��<L9N���
����ӡ�I��y�Ax��újb���.�E��J�}q��e3fek<+�{-#:��H{yq@����Vyћ���KK�A���`�6��',��� o��G�KXGlw\Y��4�7���yw����% ̎ﰀ���|MJ�}����\�H�؟Y����l���I��a�栺c��J¯^��g�|���h���L��p,�S�v{���q�ē7hA��
<lm�R�H��wa}�c�l�b��VAn^��+�}��Տ�qk�;��V��X�
`D����:���������BrVS#��;B�L�i�  �9(�:��Gl1����T������;(h�f�����	I
�u�����}�m�~~=؃t�:O��i��&��&�bkq�D����hԪ�˟�.�%�����8֪W�s��A��+T�K᥅�[���FY ��w�F�k቎C�o�IL��U ~"��S�D��wu����T�ء�^��1W@��#3�]$9�T��s�1F䇸���m���.��F���.\w��P�������1`�L��t��'��"k*m���pY�ć8�����U��0��6��=�;�]]]���$3��i)�����y�8��=vdh�q	��xI�cG�&/E�E@^������t���0;�r_1Ҧ�	�Q���ϟ/ǲ�&IL��oM�{
��L��u�7���:�+�[(���ZE��DE�W4�(��'�5�{w��}����`���:�A�`M�΢��>@U�W�G7��"�3�0|\�e	Px���gk6��5���`I+�2�~Ocg�M1+����EW���E �����ee��4���,�c�AAA��j�ƈ{��i�$O����|(�y�n�bbZz��B��Yk���{�e�w�������<ǓJK^�VK&�`�1�S�|{�Y2�Y�(�c��mV��4@p<?�֖�B�F%����cv_�!�iLP����W���$ɂ-|gML���J8T/N],�M�d7�975t��|W�<AqP�d�����,f{�n�Ch�=�W�_	�[#�^�����x��ڀ�;K&�І��胣mj�!qw����'~�dwc�7z�A��ބ��t?��	�M����@��T���y�M�����FZ����i,�����(�p �����
�`�C��'�_|(X-���uh,��Z'�?�ځ�L~t�W��o����P���)�qO��I+�(�ơ���֥�ܒ���~�����lУ�����V��+�ż�8����	2q�)�Ѣt.eQ��#gqq�y��Kz�Y�= �P�6�-��5�x��OPk�����R�>�?�X �ޚ3����*�I��h\ N��Y�������ej,UY��Ej̆�aް�?tZn��k�^����{~�Z�$�P	�'���}�f15`�j�ܯ6�!wI�,L����&ͭE@H��=B�g��3�w���[�ߏ\���I��M6
����{�H�}ë,��r
	�:�m����% �Vi�\��1m� 饤���"��1�r ��y��Y��QFzlll�VD1M��\?zT�K�������H���)���iʈ�(;h `�Pҋ���
ƹywd$Q����mO̗N�z�y�u��2�V�x��?�\��m�����װ�s��Idq��;�X�֩8+>0�u��uը��Y1����p�U���-��
�C�8��j*�j�<#��V.���_���A��i����p��~��LC��6 0O}Y��z�}*/	s�4���;�q��I�wj,�4�g7��#I[��~�4�p�c2U�������g:7hH���c��<��׭5J�:��܎�}�}k�B4�Z��N��CXX�=�8�0w=1��P:MP���Ly$Ǖ�_H�v�at��g3�|3B3}� 3nu�v����ş�n���c�����z�e�6|�E���:��q�i�������I�=�ܳ�M�?L�ݥ�4�nB����������ا�O�_4�M#כ_?���tni�I����LȄ^Y�����3s�	$�;�����̮���m9c�^}�+�����!��̏%!�`����c�@��iٷD_�k^c&l�������P�i����*`2{���!%Em���Ƿ�K��S��UO�?��^�";�����H��AB�ev� "Cw:���\���q��<�_hq���C<9o�oU�0�W/Mq���>�HϏ����B�8Xǲ๗���cθ��2���߷�Ӑ�8 ����;�.\�RVQ(r��y��-HpW#U=8�N��a�W͛�Rw,�_��NM��`��@.�����<�SK����7a���BW�l3bM]P� ��ʇ����H*�9:+��j�nma�������ќ#9�a#e���V!�HVh ��l�)��I�u�<3�h�欞��Z"�rGxz���zM��}��e�w��Ɏj��qq[����D�C�2�� CuO�Yw��=�;}�T�R��fT'M�7r0�ڍ"p��^+�O����܊�� ��ݐ1>�z=R �?�K�����(9��������~�=�� ���Z��Z58|)1ދ=�:֝�N3�y��D9B�h���K�6t��ebT�?Mw,�l��JH?ށJV�q�^g_¾
_�QW%ïW9A_�=��9���Gr��⏜ZB�q���9�)�t�q�F���:�z��]d�� _f<���xd�L���>9��a�Dg�u����9��CVV���
v���i��X���SfC��U��a�q��Q��vp'q{�\�%����`�Զkm�`�����V������,bGY+?�-Z)3�3�^�(�
To}�W���No�x-=�x! ����|P̓ӄ�H̍n����;�`����:R��9��=e՗�o��q2�܅��𧱛e�	:J{���+�Q�z�i�)G���!���Tx���v8h$;����_�ulz#m���`|v�M�B�v�d�_��w��f3�P>ii[�1�M��'���.<R,�����;8���H%�v��<���Je&��1;��Q0r@��eH��T�sZ�-0��s
��v�r�fOʾ'��C#�ʭ�Gj�$�(s@u�~KZi.��e܅�^!�f�,�W)fV�c�V���:\�a�	A�+j��G}/0��m���x���u�,���`��J�4����c�������=m���
سV�S����=�\N(M~Rom�4Ec{h �`��x��"�6�Ǥ��	v����z0O�Ȇ>xꑦ`�
wb����]�A�w"�}q���[����f:�O�o/��3>�;'G�<�ä��z�T��5��h��L���I���e�e��>�����}�����di����2�w~��/ѰA6��~�����]�!S� �������&�q��ٓ��	B5�_[[�c��N�DPa�)Mǳ�v�Q&���D�_Fp��i��$SRR)��b�yz4�J��J�(��@�f�*C���D��6w�;\{{�Q�zV���(pG!x�d��E��o�4m����>�}B�1�=<16�.�Df���#&���vRVd��h?��b{��Q*��n����C����¡��������[��N˝a�h�T6��/"5���5
�geE
������ж���~~���&*J��~W+�Ϳ��$��KѰJ�l�����9��$��ZwBr��<�����HZ�s0�G$ �p9��#"�?��� ���&+��Hl�c��G��b
±��b��Ɛ������� k�4t�����Sw�i|G�um�W-15�S��G��Bܜ
Ǵ���	�j�X���,�r��j���� �*�@���jCi���n@uo�v��"���~\	�ng߶���B�ڈs-`U��oa�18?9�܏9�W���̱�;� o����[���n�B�nV]MM����^��l�����klJ��i���3�h7��n��3��Ʒ"#��r�2еUw���z��Sl���}�'�(�<�d�j��3�{NV�p�hhdȳx=���>��zr�R������VHM&`ݣ�N�Ed�?� ��&ѥf��2,7���]U������b��	���T�%�]̷_ɕ�;�?-C6�f����u��WV�9���؜�1�{7Xk�*>,�~Q���$aq�j�\�Z���:��s��)�����X~ԯD)�k�	�-V �r�T{�4t��C��%H@X8�M������"~Qz�'C�����S�I��e��|�=�_��޶NCy�FA�b�r˗>O�e��,z�D?Eף��'L�6��C����ق��$OҐ�!V���m.��@w�G�~���B�C\��C�#,�@�LPZ����0�v�T���R�P�PճR숵�raf���{�5�e�m�u���,��`x�]�P�A�i��E5��4,ߟ	(Wq�J/=��~4m]�U.J�1�+���g.�.���**M0Z�u>�s�$՜{���v��Q|�S#��پ$L�V��"��*�q��4�c^(��~' �N��#��8�*`
���<6�|���p��n�+��7`v�>4���0����Ό��d2��lÜ1�y3{��Wc ���O����JG7��/���ן֝�BbG��a-/ŝ>��gl8��'u�N	4����~��YGYA���WQ	���H�����'��?�C�9���M�ָ+����r�,Y�n��'s�,c���;���Ii����P�R��������$/��N�>��Þ��h��b�\Jܸ>�l�?S���(hl{U�qR:$���ׄ�����/ߟ��]~.�o�u�Y��"�#m4��ۿ�JJ[�nG�;���^�HC��u��~E���?�?2��,G�$i��bnͳ²31���s1]��<��hV'Ʃٴ�1�l͙bH�;j��t���B�m�_���Z�q�O��1�����;׌9!I���Z�"%4��M�Q���m.K��>?UvJkm����9�#v�agc��[�IWCC�k[�޳z���[>���1#��xƥ�Z�2w��J�kb�Vv;����.��rxD�l��`��ዚ1�\�3OA�ZZZ���<�I�=�Ex6;%� ��娞�h�8[��+��%�
�����;s;��|n>Y�� *�VMu֚��p��8ދ_�I�7�!{ qw0���SڥN_s�I��;�����阎��w��i��g.*"ۮ����]ŏ��Ȭ,Y˺�]rv�AlU��������w	�o�d��׉*:��bM��ݡ��k<�A��U���e�j,�z�t�3M&�����Z���ߋT�N�ɲ�b��W$�RW�%?��ԼH@���|�A�Gh���py���������D
��]"˫�ulZr+���H�s�T��1�ϥ8OrM�7��%�'�5:���^�R�!�@�����{f��2�����£b��Q�2�ؙ$ҽx���g��)^�ڷ�oy-���+����Í��}�ظ��2����$9yx�cBk�p<=����m2�zp��Q4�
��}�ݲ}�Mv��o��$��;H�޺����i�W��S�����T��_���ꣁĝ���`yi�f��cONs�����Q��snL/����ͫǟ<�Os� r i���훂�������4j�e;�U���tл���ɋ�#h.�Nc���:��"�axdda]��:���n���4�uZ�V��8�"o���$4�䓡���r��KI�x��_|�{��8�aw͔S�%u����S@��@yh��a�}�?��܆�z�F������;g�8�;�b�5�� ��psn<���Yr4;�U
ܑ���g{��Wq�֨�����)_|Gl9j�FǷ�K�+�]~�|[�L��p�ߴ��ڲ(�������}��.���ut؟z�!�I��-A�	�9ո\�碣]���Y[snyYJ�<����W�a;�*��\�@/��Ų$����yO��@�O��hh��Ԍ.�<x�=���@����I�Ʌ�P��4�i����/�?�; �of/�~����³���xGkg<<#b���caa![�bE�˫�vw�hM�Լ�s���ҡ����-���R�q�C��1�3k2��@,��� ڪ�2s�=L�5�\������s��(�D�	��n��W��]��n�r#E�M}���7��ݢgԌ��:��
E)�����ɦ@���j�������Uꂀ�*,q����2S|�>y1,��Z��S�F�S"�c�4?t�\(����s�%|�S���o��e�9{Ѽ� �^�y���˧��n$(/m.�As�S}Hb~�}iq�,u��������V6Z��ܳ�k�xf�mK��aWeh�����wu�wR�If��P�Y�Y����0h\����Qw�$*���)ҰA�]c�0��%��"#��F�k�8?8%�����3�����d=����j$ԔʥRO_?A\Bb`` �Er������f&_)�L!�=��hydYHn���~�M����L�ؠ,�H%����t`�?Xb�Uu��� �ao���*��;`K�!҅�g�2��'s�sVK�r�dC[�!���V� ں�V�Z�K�H]VV����2n�K�ݵi�H|G���4[�ᶻ���oc#���>52�51GOE�kfh���2G����޿�l^u�6�ר�����I���Z��ighJ輻�5�M�;���:�Ö�g�C�vt���GJ�l�� NN�(�<��+Iv;[oΏT`������ʢ�Q5����؞d�[-9.6�\�Q���Zφ�<��������}A�����=�B?R
V]��5 � � ._U��fݧ?v�)�뀫�bԝ�216�y��A�5��ţU*$n�gn�`�����իW��� �L�R]s������4��S������^�e�z��PC���?��x��Ĭ�W�����@֧t��d��������!]	7ln�`>{vhE&r����\�c��'��8�"���xp����&$FF���K��=Е���lii�T�*��H1z��D"ָ��F�:�QW����iȹ��GETz$�X.t�l�Տ�;>�g��+��{[�m��2��A�ZZ1}G@�e���YL�p\�* �H����׿U�1��\�^���*��׏*ZV+k��/^�---}�"`���kL�4[:M��QƝ7}�����َx5����<'R���r$'���Gs����L���Օ���L�S�!S���v�_�C����ٽ���k��me����6NN�GGGׯ����y{{;���;���$��±�[�� ��a#���J��o�Xo@��Wz��**7�o��~*(,tݏL阅���>5�,f��#!���߱(��\6�"��J�3נ֦�;�X���Q.������hGG'''�S|�#"�/��P�-��h����j�c�S#��6'I��"���Յ��KE�Y��E�#]���3ϻ\u蛡� ��F���G�����������9����@��N{�Lm#���5O�_M���ڊ���o�z+��y|�<e���G,,����n\��zf������T{�6��� �o�����j��*oP�f��N�3��LÚlG'p=11���1�=��W�͙�4�a��Q.���_����P0z�{O�'f\_����
��:���\aG��K�+V6�8/�����;/}��S��N�ٙ��?X{�e���,t�g�{��"�M3 +�TT3w�S�B��-K4�@��Tn���o.�Z��	 Y]��,�I�טE\�������w�xoWd�5���s���㯞�����7Z��"�>��jGˠ~�u0Ah�k�<|�^.T}&�99O���틞���bb+c����G7�O�%^I������@A?
�/����L���7�$Q�GhM�Bگ9F�]��PhVͻ}��i
���m���1;~�������6�c����:N�=�Ј��� *
J�����}o�EU���JǉTp&��ǘ�0X#<)�}�d D:�x~��u��	 ������T[ϼ������6�BXR�;N�${�ul5�2����<���Y5Z�����Lb߉%�9ɩ�I�n7k�j����sI�+����'}�BDi�q����� �z���aRBZJD�D@Z��F)�Mw���l����DE@$6!nR�- �����|��k�sTp3�ֽ�{�̚ƽΩ6���
Q���v������Y`4������`�}h8�vw˵���y�b�����!�A��d�d�IQΝ�w�W��<�QG�rEp-ź�eIA�w�����Q���%��-����E��v2��;)��@h����/��%jY6Z�X�SW����Z��#GI���	��k��Q�v�9j��z���w�T?�W���qE٧�W�VW�n�@�F��<�)�(EI.b�S��f�A���k%[�"T����u��	������C�\�5�P��,!
�$����ö�|&���R�>��m�E�+�&S�ʕ��ҷۘ�	�2�<�dx��gp�R��oVW_�a(�a�䗾>6^��y��D!|�!�]��iC�'��f�5U
�6X��좏����Rj�q3s�����;Wάx�%Oj�2x�S�M6��������K1ҟ�73�j� �[�'�����tM�"*TZv�K� �m 8���\R����5j�(r���A.��MjР�eM_w�v�*y�p�\��"c���M�5�����g��+,++S�=�O�S�1��T��d��]Ac9Ӏ)d99�_>݋ �d��$�0GX|J�%��f�kuI�R���s��op�ۼ�6�֝�1��Kb��갦553����˪�U+���ګ];��hZA�����^(K ��r���E���2����X�^k�}��WcQ;�)w=�P�:��J�!�u�3�fNR��.�vnߍ��}Ĩ��#^��=����Էc.�!��X���)�و�n����u��+vŬ�hڝ�R3$��G��Yӥ��6�����Ư�����g��v��8͊��Zo?�a��*D
�B�+�*T�z�EĲc;�R^n?U�`͔�h��@�kG�$q�ɓ��N ��K�@��Y��<��@��ڐ��-�I�a�r����s�s"��[�a��Z���;�T����+���gR˭,F9�w��x�~r˃Y�t�pB���l����~�:��p��/K���*�=G�vM���D�][L���r@tf��y��%I1R����`!�7���֗0o������T J�{v� dle '��kl\.O�k�E5[�t ��ۨ�ˉ��z��>(�>���ш�����������&�TT���*��Z[���d5??�$��t�p!��epӊ:�/�ֱCb���[���[ќ������r����Yf��g�~'��ss��*O  -�0�:+�<��Z��^�oOOr|���z��;0%�m�����|��T���ד�/���d`�`�|gyhUQ��AHD�
����{_X��<����|��M�i��Hz1@0'���I��~���-6����0(�:����ݲf�1��'`�x_�3�%#��D 3%����ˬaي�~�i���F@m%ɎC�;R���p^�Z�!@{g�)Lbq��)�J����c�R "�s�V��C��0Ϫ�m	b�/�@�@�@�Y��n@P5�.��cT� l'�>�4�k��'�W]�v�(���C�uT�j���h�ܱ���ぐ���S�����!�:W��������Ӡۻ�V	;��I?;����5��~q�J��"S��~󴰑�A����P�~E�����o4P| ��=��m�N�ΐ�q��=8�V�S��k��ؿ�зl���v*�j5n�#T�ǩBW��Řg�Vpp`m{���k�'��ME�}��.�|��|�w؍Ilu�s�䭏x�#o���:�]�_��'l,�
�M#cɺ�+mv��+2&FA�0���v�jh�@�14�]������U��"�ⅆ�0�q�<�oS����|��cg��B����	D���w�/�aW��������
�#��-�aZ��45����O88y?��8wnj@�q�؛�" �{V�{^�N���n�~�`�<���^N]kkk��N!���x����}��R��<<t�g�����jqlJJr���о�Z�x+2���n���eIq�
D�� E�c�3NM��fWW��;v|l� �Kߦ����u�(�nX˖�o���CJ�R�XY�2�N�o<|����Ttё 3�����@3��� �c�UH��|�MI�#Tc�-�f��#w������1�NV������I����s�Ͷ�U��ᇏ��Yy7(�M̩?��a�*�3�I��O~S-dz˨���J�)WK����
T��}�"�����A��s9jק��4�vIC@�ʁ�SZ\���L׮Q��H��j́����+4��g~˼�\�m�1�Vju50c���93��EP)'o''7>���J�2@Aن�[� JE��~�s�����ݫA�8�o9>:��=]�o�+��l?]��10� ��* P'�ù�Ӑ�W��ȍd���k�8~��P��Ic�����r��G���}[Z�b/��P
�� 9��;9i~^�N�Z�Ĉ��������>Hao����	��ۃ�Ji��Y2	=XW�wþV��q�L|)kS�L~�����9M���pWS�܃:���.��+� ��n��$�8���$�5�`������څ����Jok�
���'8g�w:T�?�Π˝�%j���4���N���F%�:a���ܬ���[^�n8|0O//��(����:(��5N2���3@h�H�;�*����:���a[��s0��Q�GÄ%OφF��g�J����? ����kV��K,��Y � l��	,�o���a816ZqѴ����v���)t�*
ID�hX��j�S�AK݃r���b���n�A���1�+����7@�4����yH�<X{���z���0�g����'rr�P�H������P���vv��߂ ��?_�Fz}��ȻH(3�'�d dñ1m����x��*���Y@�Ђfn�s��ppk�� Q�5�s�����KK�lɴ��׋*U��28S��D��%A��#���~�f�?~���w� ށ������!A��=T�
0�
��8��۞_�/�<7%:��IgC���6�Ɋ�'�x�2^T=ym>��r<::z۴�b���g�e���貇h�j�P����g��KH� ��RU�x��q� ~Z����M�c�
cۜ�+�υp�Gt���6>1V�j}��.}�]=a�I����Uo+���P���qPa :��1+&�~~���PJz��]]ݹ�O3ϑ���箇V��:�����w�! �K>��m^�JVRb1��llo7Yt���6��#�2X;>2���N�|���v�3�Q�[ݴ��Ő��k������H�B=�5eF{cZ�7f~'�b���Vg�^��[��)�/�{��[�'�m7^�[
�JP��<�Df���4j�lt��Ҿ�N�jg��D=�5��>���?��8�bX
X��_����C��b}������ �$k9����l�� W�B��j|_��)~��Q�����Y�ÄG��o�]��-Sa{���&�}X!־��KÕ�vxv�1�3�ԭCo�Q�[Q����Q�L���֏&TM��eٹr#�)0�~�~S����TV��2t��
�h�n�SqB���\TTJ� ���-Jj՜��.����-�C�4�7��D����"K�(����ר7n���X��-�OІm�����@�\\�A�����ly���� M��p��yoooh#U��)�lm(@�
.���t�
���
C�(��2��RΘ��Es�0H:׳��R����03\�]��Ó?>T����: ����3#ğHB�����G����-�k��TkkZ.㣐�AK�W1� ������oCű�'�9;�>&p���:70Ѽ�ϵ��l�u�B7t��I����ڟGx��p�J�:��%x����7��d|�	@�;ЫЎ@�I�K���EfV���I��;a����k�*����. ��������&�(���.w����*� n�pvgk��4G���wS�n��Uᜉ���241Q11�=�
�a,t��p�������&��H�AT�SκIL�]b�c��O2�s.��������H�4�{p��w_�������=?1997��' ��i?�4W���o��Z�%�H��#�?`�jy�<��+P����JaL
��[��*���ӵ��S��Nש���3_�?z��a'��������Rr}����tvwM��mhh�Ʉkk�������yM�1.�L��ӆ.��w�D���R�؍�+�m����%���'P ��6<C�끉}W���з�"��@SS3:]�w͖V�F ����!�XP?��j*��9�΍�c~L>�����m޺�3��ʻ��Z�9�o���_&�-�6+)+O��'���744uudffg8%l@����Q��ķ�6:���WD�\��ep�����6��P�V��R�3T߭��X���y����:Z���a)����5fL���0����8�&�^%̂��
m�9$>��cs?R{�s��V��ON;�����)��@��zQ���)����iv�Pi�2���c���ITT�9��옘�����������c�������l|z?Խ�qYRH���= 2�m�x:1 V�o�PC��$h����u���Z�� E�d�_������񝝽׸��'^�m`�:i��u���h~�t�C�L�?���։?��i�-�~�+�(�~E�JY1��VO���t)��/m׷�&��P`�ꉵ�@��_.�F��r� �.}ئ��o�%�@��@�yk�N:�k��]y�C��������k��0dB|k�6e&��~7sM�����N9 �|9�q�2��ep�ˤl�����w��b?�5.�S�*@\���_�hR3�T�����[L7?������r�pw��D|�����S6?1Qt?pCy���M��|�I��X�f*p3��o���'���1����.p������]��	�'u�ܱ�����3�Y_o��Hl��c9�Ċ��|q�A:��Ί��]���c�{�`rS�P�SMr��ȋ��,ǋ�Ϡ�H�V�!�U �omm������p����:A/���d�y���Q�F6o��`*���ｑ�(�X���dn���������9�}Z�,P`Q��
�� �;��7F�������B<ζ��SRRn�(�������c��%;���ڀ��Vș��Y���6�p��oRp�>Z�@D/���a�kV�frV�;w8ZעWƠ���<f��y��cb�=6��W}Q�M?,8�h�HB�$u:6��3��_x�*���ԤT�6��9��A0���]*�`�T��h�����@�3�r�@�ж(\�f�̪]�!N�bv?�I4���5_���=����v�T�.-��s��1����9?T:
�Wl���5D��k�^Cc#�U���Ufqfff=��fM?�Rg���#�~��lvՎ��՟���t+/��:��G|�o�[���!b'k9}�=�eU=c��j��Jq�c�X������OLOg
552�1�����=$*���K�$���Q�K���)޴�՘/I��sT/:UNUxz$�?�377E�B7��VsTVX��l�jG�������g���sq����[[Em3�sB����:&��7���Q�9�C�@C�p�j9:>V�C����}��h�X`Qf��c����<��Q������ă���\'�4&���������x���ٽ�1��h6�w�ޔ��g~�����߳VU���7w
E\�5اlnn�O��h���@Y�C�Tyi�F<��}�ZY999�l�G���O"��%�+�F�摥cG���T��J~��YBozf<��Ϙ�y���3�qkL��烦��خ������2l��oSxW�f��������LYV����V�%C{���s��s-E{���A+햷�8��s���S�U��3��������+����%�
�''g�R���үb�%���:�f���W#��[NMƃi��z^�8�M�CM����S}��FyAΞ�9�@�|ms`9�ҿ�-8V�^t���Zƽ��Z�K�΀�9Ѐ]9�I���'}+�g֙ŀ���+�f��|_q���*ooG�Z	�..."��\�d��%�3�{�z\-���yҜIݰ��6��$��g�G]���iT� >�n��5����� �yG�I�߿�<�Q��q��z~

=����i�j����7����Zo 9��L��n�_�o?�ӥ
e�Q�?�z0I�G�/��������eGkk+�i�Q�ؒ�їC�[�}K{�4 ,��/�ЦU.H��^gr�{���c�����=�M�T9M�3�ͤf���t����M�7\��j�}5�����a�䰵�uYU�V��
=M�T^~b*�b�6z���/W�gA�y�;��`�'��4z���i��Fa�D����z����˹
��1C������,-����Jf�(��"- )7Vc�����[;�g�g����:�lub!ߣV$ظ�0�z�{��-��&�9'���ΒQ24J�yZt�>��12���;cE���2F�V� @n��Y=	�|($TVS�yu��ЕE�[��ϙ򦁥�:(S[[[�_H�ek[��@��\(&���[��@�Kl凜]wou��!��i�<��w��\vB6B�xn@'��HB����^������b���aV�Uz{�C(�\9���KU��
��+���u��j�|0+�.q/���B�k9�����:݉�!��ϼ��Fr���@���wa���u�a�m~vw���
:ϵc���F<{_P CAA��� �z�8�)h`J�uZ����p2@���u�+ukM[��<�6V���UX��=�J�?�<�)�M�ϟ��@�&����r|���Q�K>�-�i\�B.�"����$�=�	�^~��Dl���,^,�Ie���}��f�|�V\�	�c0��گi���ܦϋ��KoԸ�;�~�Gi^��~�|��Xс;�8 ���Q��� I�Ф9�^>֘���>h��P��ܝ�����F��U�p4��cL���Qٯ_�b�KU�7(����By�:�T2�s�p蛜�w�?����Er=�)3@oAiv�w��D�c@�{n����������x0j�eH�4@��ԋ�ܜYx��묟�ƫ�R�F=c��;D���r	��t6���j-;�q����oҢ����4ϣ�a��U�۹�cS�`Ri�ݗ���� �)|�R��~-W�n�5����(��峺�v���s�%k�"#cc��k\B�l��s.�l�c�8Y��u*�P��.~69�[�U�~S����9�V�d)iiPf ��;*��l�A�//%��-�	��ß���T6�A5K%v���6P����A���ZU焻R.���`�w��^��1��!%�c:9��C�	���CE�T\��rA��ކ�5%�Q2�������vߣ8�?X�`t��*��~���dT|��s���
�CpnJ�bod����z�D���4��$BMB�
�O��S�UM��ߺ��Dn��p�z���籢~pj���K^�NqT��z�	)ݲ�����.z�Ey�辜4˕�k�x�5a����5zU1�$�=<t������XR�L ����̲6ϊ����蟼?G&�WK@IFūA���b�&��F��*��\�m~��~��xQ��-w�o ����ٿ��V���v}Lļ~�w��v;kț����o�:Ď��e�5��@B�7"Q/�h�J3�["�Y��M.��_L�ݮ*u��@6{hp��Td��_�D�Ȕ�ۇ=�������⟘ӟ�*�\"l���J4��a>�ք��mU��G[HaM�j	*�ѽ��_�����34�̪�ǰY��Vm]gb�tk�6� 5��?�_�]�'��^���d-����T���L1wO��Re�.�T�p�K��Wm�;���~��GNp�f2I�����v�t����ᗁ�v���~u������ÒH�ƃ'DE�ָ�%�P]�j��0L�1��~��D7�J�4�y}^rU�wf�}跲�c������˷���z1��\Ͱ=��	�A���BϫV�]F���e�}��m2���-���kcb�V�%���0��3�(�m�4������i��#yM�Pz�������԰0����kվ�*=�j�P���sv98�#�<��O)mW�w]v�G��5��=�\�7�%����<;ޙ�@�4x���C�c��� ڵJ�{KC3����38�B5�rļ9�v�Mf���I�f@Z��k����*��8*��d������1��r*5��0tJ"pbzU�8##��㳛�ț}|��e�w>���@y�?]��/J��Vx~������[[�|�〭A�^��`-/�l�}?�>�@����4��J�߉a�7�#W�ԃ� d�*�V���P�by�~ˈ��~��[%����ܐ�7�z�aA;݌�Ig�W��j��6�ʰ�Ȍf���Ub�gvB)��,]��-h{{n^�!m�ʔ���6����������+��&�K��m��J���K���3��_� �֐���qj�l��9�߈�J��S�����Br��V\����@����i�o	R�����1�{h@�C���������V���gn�E��ۋ�r��_�SǾҸ8���,\�A�}a�W�ȴ����u$йPa49��;�w�)P[�j�4V�;��=�vC�83�d�X$�t��4�m� ���''�

*���JUq�����7�;�����E���n(��n+&I�#0۩~�����>G?�VH�qO����>�
1�?�ׁ�K�R�iv<|"��4�ka"�8��z1&6Q�(EI� K\h(�
�O�GԒ�V�t���K�wrw��z�TIݶ7�ᨋJ��O��Nl�yLOm���w@�x|b��r p�&Wb��4A��0���q�ʕ6�2X�����t���@jL@Hkjj����V3����ѱ�O&�.�(�Ǯ"f��t%"�ľӊZ	�?'�b=�3����+�3G!ۼ�ڭ�Ɏ�S�c���1m�Pxm��cgg�5Lw}%~
���}f��Ѧ�;����iU[�Y���v����?A`p����C��;8L��U0��ƮC�rzz魭-xU�_��}9�o� ����2u �B���h�k�x�����`�D�//�5G�{���bR�XG�)��i��p�f� ��F�����*w2_��ZUg�8�Z��� owv�~]s�����G�EZP
�����&D_	���϶^��R�;���?A��7�|_��Q��<����Q���W�cp˻}��w�Ӛ���@R\#������ ��C��(��zc�||v�z��C��R���7�T��z�1_C��^����7wϯe��3N���[��w5Zι��Ҋ�A6���(��<����{�H
�&�7��:��O�/XR��� ���ŋ��A��&Y��?�҂<�7ea�>jr�i.�� T.b���O��q���y���4#$$,���pa� ������<)��ќ�o�m˞�6d�ui����R�xM�~�@+���%��"���t�>�V�/�lŗ���Lڶ���n���]�R�y�g;kj;n:�E�c�Ꮵ;O�Sé*��ٕ�|��k��t2n�sH��Y�W�tݔCf����.ccTž8�#%
���u����x�k�μ���Ey�O�_w��կ�Pl��;J"x���[(��6ǳ���?�r7���'g����ߘ��m�93���L�-;�؆�ӧOߨ�zušZ���)_��bzܝ�r("	c�-�#�W���sg{��^9�Zv��-RRRBF5��XkC#�����j9�����F�P*1[*���bS_��0�ޠ@�m����L��fr ljjj��g��uj��&�������c��lpn������_Q܃g��Ni�d�T���j}֓sC� ������k��S=O{��"O��P�msZ-�H;��n�1o�)o�I�53^ll,C�
#9>���e&�RY�gƲ��{7%ɲ�PK:��t�J)���uT+�h�OM���AC��U�~��m�������kW��֖_@ ��/��#�O�/E�\E���:&H(��\��>I,��UQ���Y��Ls(�=��J�R�������i�\�M�Y�~��e���A��~�t�6�!%�L鎂��vz��g�m�u��mCرv��T�`��2m��`�5۾�+��1P0�1��� ~O�f�C�+�*�H����V�n5+"�a�e��F�+z��]�ӹ0�X�Q˾�@`wA��n�Tc�͉�!��-�ҕz� aI�\O�������Q��ks�\$�T����b�<=��ʺ���~r�/Mŝ�bV̉��n�ڢ�ĳ��Ӷ�y�ć���?-�Ҿ���W�.p'|�{�;xCt"�$L��r�<ԋ�~��\��N�~��hy]�g��A}���o�����a�s�3�n%2b4x���7Zg�665�ttZ���O�#}���(���/��R�f�!h�~t[^g=B��d�'��_ؾ�L*�}>Y����0~�┑9���X�YE*�KO���-�_��UFK���������pS�"����204�98��Y1i��q�vh��Ko2%�<��=�An=�� 1�˖�i��f���0l"C��]F��:�g���9�К�>{�7�$~�	cA!i�e�<iT�i0�p�!�I�pO�Q��x%�'�2k���զ��$�R�YxVz�����
BV2O^��PS��Y4Mp�T��7�q�{�,�od��fTIiT9�$�-م�A�v�mUeˋ,��^��`ꏞ�����.{�`NF%������y���z��o�1]��#��"����9IhB�»S�S
�I>�%�u��A+���9��f���2O^��˻ h0��V�nX<�D���o�
�Ka^�ċ1����>I�{WX)�ݬ=�]���^z��O�w��}���q��!o�fƵ���b�"�τ!��ymy�-���� >�*�W�X9r��e�����\E�i�\-)�_|����>������=�5����ig2�z/���:�1��+O~la57E{�JT�]�sX�/ ������:�>W�vW����Mے��
�`V�<'.��������Kw�����m��&��xF��2��J�zJ���]N���N-@��0�����|?���#ؗ.ELp��;O5e5�[�Z.���".:�I�
��:<=�{G��:��p7#��`>[צ�X�_h<��˲k;��RG�x&.pA�]�U䎽�Ӫ�������c_'����M뼊dV�s(ܼ���(��f�a�>�Jmd�Ã�!}��m&�t�	�ӷO���e��'�uu'���,��������f�b�_T]'�A���@��l���I]N��x�y�'���
gN�u�����wI[^^�o杻���ΐ��v�>��j�VY㘭���=��c�Yu��nAU��C��.Ů-��[�n���K3��Z���0d���E���M�>�/��T�ݐ+�#���DKg=)��ʱ���00���ĥ!��km��8�m��=�B���^h��=�}������)�ﺦ��e>��M�T�4��x�H�_X���#�=1|����?yZ���H˂9ʲ��.*b���z�H[[[��
��0A����0Ѹ���>�ّFˢM�u�n�F6�����w
��,F� q�ɻӁ�C~���13c�,b[!{�|
���~�]���Җ������)ACG�zZ������o���b�Aھ�uӲ��҅��=QQ�M\���G2_�hlo#7|%v�]Ò'�{f���Zt�I��L�����p/DW�V��E٠���ǟi,[`�;��<�i�#ɚÝtg�����i��b�O'��6C�����Vr�ӣj�-�H����R��Y[c� ��:������J���������Ғ܏�_S�Y/ϖn����V�)fWZkpg�������ݶŶ���  ����<q	}_s����
�tɨV���)J�'��|�{�9Ue�(	.���8G�d �)f�?��� هl�v����{r�`�Y쮖K�x!��H���Q<p����%���ka��)������;-��C��M�^t�|�� ��G3��aJ�&��b��H��j����p���3nv�7���$��г}�l�5or(��6��_`X"�B=ww�ellL}�v��23���Y����c��O+�i�@z^�}�ЫĿE����-ڀ?=8/i��nɼ5�tww�g�.�$t���cCKC�� P�"�R�9�Q�G[��I�^�z�Sqzyq�H�ENqߔ��(�Θ�Z�V*����(�\�ş$U��-!k�����ڑ�d����7�.*����X)��+�4̜�j/Q�
� ��ҏ�Ҳ$?�ׇ�0;5��M�ԛ�`��'���V�R�-љGeT�+[p{BlU}Rчe��m��n|�H^��J��O}S^�(��O�\vZ�����I��r#�֣p��i�6��ٿ�C��?qJ7)�{X���y��}�����*�=˕��n�w��H�84ivA��x_�d�=�rH�g�4���j�!4iqþ|�/$$t4��Ԧw�I�݂w�6��D=N�Wf�?9q�����x�/��5��2~ϓ"VE��󇎎j&Z���������j
�6ۻ���.q.LFd�2a��Z|���_��
p,�Q�Rt{�Z��w���{r<cn̸~&gܼ�[�Ўݏ���S۶w��%?z�	J��[_�q�_��d�h[c\T�y�q�`a�T���)
��!�x81e����B�|>��an��#�-�#�z���pU�ez=Fا_�m�ުZCwAw���r|�Iد yȑ6[I|��c�>ߎ��}G���n�3j��zOOE�J�Y���J�U=/�4���A��|�b����>%=n�������RVVnv[��2����d�.Ցʒk1Y�R���3�#��(�^z	1x���,a�J��x7v@v���$�.�2��}��M ؅��
EZ@sI�O�1nZ{o'�ƿZu�n�E��@B/��mX4�E���X���c���ؤ�� yY΀#i�,'����4��|�$�Ik��1b2BsW�HR�
4�5��Y��a����٦�5�"	�}/�H>fA?�H^�\��l;tz���?�6�u8�������p�gMz̚ԣ|�#��v�-���{b������������~p4��yUj�{�^��x��;9;���9�
�H3����ē������Y ���O��>y��	:R�����tz��YͰR5��K__�
k�ͨ��E���~�V�]�	ь_p���,�LT�@�t�m�B�*n�I��0���-Mw�88��q���Q�V���Q�^7���<��Jw��v�������P�?}ɋ�in�e� Ģ�"�05�U+�۟�����=�� �FC[h�MMM�P_�%��=�H�t�P����`t=6km#y9�@��o
צf��T4�KWQ]��ӐU-� ����b%j��B¹��[�Ehq�bTX1���� t���sIO�kҝ�.��� Q�OJ*|�	/N��v��M#���bE@P��j���i�Ċ��{�z��M-6J���Ñ�8���F+3���i9�ݺBL���������M%�o��%`��wc�}6:n�����e�Fm�`G��0�e��ý=�_�>%����Ҟy�R�~����$�Y���ݾ�5hn��m?���q<ck?[����������9
0�e���cwZ�p������X��1/]�>�$CL�8���w�4��K���3�ݕ����S���2�����#Tsgc;F�N�-MP*=�R���S�hr�ѫ?B���ho�5h���Y�1ߵ�ӥE�'Ѝ�h}�[?e���#�@K<�H��S�.����g��~�w�l�4H�[	Dd����ѝ�x�qy�JF	������4���w�f��o"��4��J��v-�5w|��mN� �� ������{Z8z�̽�a�������E����R� }��=�qooO���N܍��»��l��K	RDh r���Ax����-.jݩu��_�Z�fIF��w\�u�+9ő�4�wo��D�����T��]K����F�+־���4r$���T����L�f�z��~�bbܦ�] ����p���qC�ZbACMU3�(��Qc������F�%�i�i��~�◔�`���ˋ�0ͳ����Y������;��A{��kǙ�;˧��`����E)�jA�J���,wq�j�k��t7p�3��)RA���V���'E���6	�g;]	�KPa#�	������*+m��#R͝�F��U.HU�2a���F ��47�G߈ ���;y���Vm�woe�m��4ޏFS0"���~�ES�<¶jSS�k��Ѯ«��)������9(2���$��`i��}'_q���M����"wp���ʟ���hoTX�����|��J_������l[���~������ ��M�Շ��P�|���B�C?:�ٟ��V��/9eq>.�-���ͤ@F�+��wz�:�P�����9�y.�L�S�]>��0u/:�o���R��� �p&̞��.�r͕�a��l���u�)<ok�G�Q|��]ϙTzQ8�w�=_D�A����.c�呋�P����a��t��y�Yr�L�q��L���/_nX>����3���L�0ē��4��*K/��:55F�� ����m�Y3�.��&�;&D�|��������s��',ͱ�5!���j������������^]~c?�/j=Ԫ����^o0uR�Ļq��5?��J3�p���\���~Xo�l���M�R��Dl�GX��#��q�܉�g)��pzG

5
�jy�v��a�3
�5r$���i���vO���H��b�JF�e�>�����X��~��ٶ�}K��4��c�9���CԔ����wQ�)@#66� �<�MJJҘh�Im6G8>��Z�Am|{�*1��6+9ײ���F�^��ZMK�u 
����=�S����~�;	]�G���﯑��Aሔ.��*vr� ���@���<a��0�(����~>?w�k��'%�?*Xͪ>}��gAp��޷��#8n�h��z�$�/�5��������S��۲�L�#dI���.e�p{^Ua)���y��#��4;x���㛃>�]�m�?��@���*����O�11�7A��k٨�&���YZZ���ׯ�@����;���5w���5��VcdO���Nf=o�4������p��7�/��7�m��Ode��UF�(a�h�=�2a�~�<p[���r�|�*�������.�]O�t��Ԯ#�q��rȤ�0��0�Q��/O�ʋL䬣XP�/`|�J�g1�����90�7G;!P N�����#%N7�-�{P&_c�\��p�|β��1�e�Bg_K�k@*@S��k5k�bJT����"+�����-xp�rW0K�q�� �'E���Z����ڑ��S��࿋�3����A
0/�gN6
�s�~�ʇ� �T�+e��yX�=:���&���C{+9)a�&ME��A�p� ��@,�����#a�	~����^"�����0�b]��$5�t�I�q^�����ˑ_�4,�@��q&�{L�����1{yNp�"-���R,�4��^e�ؕ��("�u8pv��0E����ɗ@v�n���y��f?�$W��7x��-��(n6�z�ߴ�ϭ�܄!�[����l�C�ڒ��[^�Y��G<9�:g 3jk�cT��d%��X3�m��M]Pߺ/���d�����9b^���[QU���w��4��	��r�X|B؛�L�]*4A��.�)��W��=U+o#nǸ�?z�)��4�������S�p�ga�z� �ג�%�:Q~o �j���s �,�f�"D�4����p��S�a��dI�l���N���6�~4v��+i���l�ͱ�d;:��jB��0�P��h�6�D�ڌ�ӱ��z7Ě`#�y�j:;��c;���9EU/	-	K��k��91��9u� Q�0�q7@�	E��?&`�ilaD�%��2����[��H�)g�铙��Kǽ[��t)C�ϗ��S�c�d�����ƞ\aw��*����K�s�.����]�a�����	�	����9�u1=-��O �H��2v�_���F#S�	c�[��%T."#�2�v�{:߿��syq�;���9	�[EU���eo���,�����\X�I4��x_�K�Ձ���	�my�Y5B��XY��x�qw6?8�C8�=uF �����j���|_C���_a��D�S�Σ���E�7�r�|��rn�㜻�?a�g�)��E�]��2NAUw[����������3�WӦ���W�檛}�G�mr��7���p��2��mghy5E[	� 5%�!"��}��]�bͫ�.<�}S�5�����-���M:ڿ!�q14�&��
�"�S'UG�.��zwl�n��a�<$d!?#����Y����`z�5����E�����O�j������)���=|S�O{��v��Q������0��u\`�a���/1ȓ�F�y��J����O�rް:E���&�{*�bee���A��窷�B=����6��� ��-����0˥n�-�������Ĩ��KMF?8�C!��S�^�~�Ǒ	L�����둙5�l�l��(��[�M?3Og���[�l��~�wr/F?���D��\M�\,�i�<yZ�=�- �m]�{���p5L嗐:ޔ�ì��88ǘ�ࢧ�*1�%2$��夁S���kl%K:rjqZ�#=�[3`��_VD���ԡ7A|u�����#��Qү�o�]!?YO=��LH���R�7\�3���s��,I��ȕ	N����u���Fo'^��:'����miȎY�?�A�Hݜ
E:���/����q8y��K��.�iW�8C��5�������Wܼ������W��_�x�vǹ���.��ȟ
ʊ�7�F�/s�����\�A�_��V�/�8)c�c�%<��}��@s�S�_����?�aA�T��w��j�X�����9o��>���h3�r|O�Ry󟼳݅��j��x��KF�*�1���n�I,ݿC"�w�jM��KL��1k裠j�%A��| Ճpo���dbbz?a��{��d
'Mu�:�v=-����y�Up���Be���_ǡ��Q�X;gPԐq��9}�t���N1��qȣg@��#�� �E������Zn��=4L�G�z��9z�R;U/"��"=���	��(wFg� ��X�mX|_�6�{��B} #��y���������G�0�cX��p/���Oռ�iܩP�oݥT$����� X�!+�+����qj�4����������1���8�jÚ0�,_"�R���K������^�b�Y'u�6g���d�
+������p��}�Ju�� 'g��+}q����57w�9��(��)!�}/gE��,@�Wa�M��9�(�h����
����mA��PB��.IA:EJ��;	�Nii�.�����f����{ν߿��yD�k���;��c���n�P�V���j|�f�Q�3o��[��n�5Q��)���R��fM.|��=`H��nŘ�t"���4 ��*�|�G��Ls,�>�݋[�7��GQ���*��*�tO�Տ
����|D���K��9/��/�?�`;Ra�'.�P�ޗ�D���iJ�p}������c�_J���-��rw-���sn�T*��z|�[��}9cj����OP�ж繋�Uo�:�8�A��y�İP_)�,"	I]3��4d+�����nA�D�G��X�`tr�����_f��~ڔIs����BY(u�t,�%��Z��m*-�-)�Z~|~ך�H9������U��9�,E>��r8K)>�l��H��Gt�=�L(?!&)�����+P9Ej��,�����tZwF���^��B����A|��P�r��G�����Nd�n}��B�l%֒c߬�;鈙jqFҎ_FOA�E~��cR��x*�~�2b�nt��@�	�N��ӻ���k���X�
zlu�goh�V�A��I����{|e������Ajʾ�D�A�~D3���+M�E�3S����AO���m%�Zƹ����y�U$���ʋ���/7^�"��5 \�!:�*v�C� # �����;�*{V�;��%z�<�i����{�F��0&����E��'KQ"�����r'��1�'^����T���!"�6F����bxg��h�ɿ<Q�9��:�����J��%��X���̋�̋
ĩx���m|i\�G9�+9����ɪ�b�5߬�����OD@_��YJ�1�7��!�W?L�Nի:k	�g"�S�Ey,X7�֝�-�Z�g��;��1)+18��QP�q�^�+��j�\���w��P�O��5�����^��!m;�/,,��N�Y.#]:+'�<�g���I��7eQ�o���������,�0���R��l��`���Y*�F��e���󓮷��Ϲ�;o����p	m�u΍�8�#h�v&8)�����rB��Q��dkR��Sw�D�b������|�jM�Oj:!+�{F�����]��uv�f�_���ʨ��$�`S{d������#�v��X?LF�2�y^�z]�	(����ῂ�-NN$3�S]=}N%V���x� r�h��sN�4p3?h|��P��0恡����!�H�!��K���$�i
�ܝ��]����	�WfL��L�2]�9��=%�R�Z0>)#�R�S��䈼�{П��Bo]%u�Ͱ����8���wS�
��r���(���e$���p'�4oBV�/�X�6̼����{�>���`����6�3��M.���y_Jo�?-TB�1`F}����w�=~�|\q�9�&��B�B�HK�y����w��,>�Ǐ���irˏ{�}��[I���h�ŗ��~P�ex��"�]�����{|}�z]h��55E�o-Z�o�[����C�nP ʫ���Mȣ?iqpz��z��f���hJ�a*r}ٝ��@o���W����r�6m����9
+��)�$c+Ϡٟ�4�5�Va}Bq"��E$��Ե�&jf`�u�;���6ǌ#�SE��v��������l���]J�ٓ���hs^�]ى�Vz��Jd�N:�#�Z�GR�@�Z7�q�}K���������-U�bQz��$>���yK`\=�|w!��?��[/�(������E��S-��H����q���M�.�[Jl��yq�g�m^�xw��rr�l�B)�Q���鞢�ڬY���7?��H}c�U�.�n7ts�%�{з�[���J����b������i~��=�?�ٍ���'�"h�9�����m_�?o�񛴚�tR5�ҼY�i'Y�T��[-a�G�}�{�CN4�y�	��^���0���CAz�l�з[�q�����M�j�0�\䲋�-r1�܁3I�᧔�f�ժg����Ab����x�OH!8~��|�B���Rj]&\>w8ؠ�g��t��L��ֲ�6-����ѦxiQ��o��˺oM��Y#Qb7H�f��y����Ӕ~�k`���&��F�^6���:����#�C� ��- �\T��u��66e�Jq_���|�cT~g_0��}>L�e�*sX�m-4.k%�!����V�f7�l}���	f�ͨqy�����������R�g-�L���d_���˖���|R ��zw#� �y��Qv��]/߅�q�M*'�S����W�d���F�*��_�А.�ݘ��}aƻ6n;}H�����1∯A:@Aam�<́�&�{;tXd�%��s�����{�ƹa���9��X�4�cr�+��e�~�@Zc��ZL�鼝P����}q��;%*5��\:��'�4��*����J�����mٹ�� �t�i=t�_B��*����L����$�����O]q���! !�*$��{�qu�H��&B�sU���|�����V�1���*�l�I܏���_�����zC���S9x��I�����3`�Jy ��V�~ŜL\x���껵�sQF�>���
�P� ��["��i�H@�:@��� ���ok�M�[cߺ	F^(����5��Y�?��D�mlI_�joOw|dܭ��yY��A�[9�nC~�=��R�,��b�rcIf��##8999o4���n�^��o��~��-r3��B�|r;LZ�ݾ�8x[� #��1�#Q���t�*e�_�7��D��Vm9ݽY�'�C�g��+�wǟ�`W��0�o�NTy��s�7jp��`ﭷ��ك�򞅄�9]���b���f�����"[��y�f��ܭ�&{<�J�� ��Z�>�+3�,<!	���ߐL�<=͗?��� b����kk�%�ߩY�(�[���6(��^z��Ͽ<#�G����|�Ԝc�?�������Q���f�?{�6L���ð��
�G�D>��+�Lh�n��ў����֜�s���<�����������0�%>g��V��g�FFjot�`޿�����bB#ꓺ��1y��v1���)?�7x�yx�L�:���������#MM͟�~��L��"�jHd��]P���32Ύbb��>��Dj��֜A$�[j���>|��ya���]�
WW�.���O�s�|��i���QZ���L%�_���\'�*1�7*F�vu�͊:��o���`X�+]#>)�ml���s��X�ak�
��Uצ��T��_g��Fc8-_R����8ߘ3<Os���0�K��_�
6��4���]~+]�hh	oO=���9��G�}�A�n��d5$fܲ�����s��e~���I��-�a�^L��ubb�>�@�/����.$��پ1z����^�����0�!���'��\�x�n�h��x�u��O�ש~m�Zu��gл����&bA/�%�n���ޛn�u������x�� �K#�{W��~��9�� ��)j^��P��^fz�Q� �t`����b�d�$��]�����Ꝁ(��[cI=�>�>�`È���-�\�5�j�u�&�h�߫�y�.�R�������1��0�O~�?�vUa�ɢ�}�l����П|��5$�Y���ǩ���Z����a���l7�Wmyll�1��u���Ʉl&8
/J�B
��K�Z�N
���ОM1�C��8=�N���*�*e@1'66����L~����'����v�d��J��<�9�)�OR�F.�/$��&�2>CF��ZU��;���W�]GE1,��ג�����Vc@qJՍ�i�H��|*�����;ґ�F-6��27���$	�Z_<���r8o�=���L|����)|�O��F���f�ל9��Ny6[^^�ފ%�5)?�իW- ]c��ic�]u�^}�j��9�+�|�	~�E�_A��o�,)�M������'$�N�|9e���C
'�Ϙ:6�V���ԏ3�~Nj�z�Pj>2�'�����5�ϳk��WR�}3��++��J oD�;J���A�+�$�S����
ȗ�ΆJ��û��̓�>Zك[Q�)F�o�ghk{�fl�_�␑��A1��?��)�sl�� nˇD%��Rk��ʒ�͚=���%;�O�.7�D�\Z���A��Cg��q�Z�����̎;��^�_v���~5��n?�����tHuq�s-����2��bTxVkͯ�fه���5���4���ȷ��GR�(�+;�ʕ��(D��1J=��ǲ�g�U�9�.Pl���?$*/�ǆN�~Wk��fY�>��.:����^��F�_Ϭ��Y]�85� W���η�8 \I�,'�Ő#_��j��r��C��-�}����a�=����/F~��Sf�$�~/�y�����; %R��D�qӝ�k�����U��PO�Lb��p�{�wB�J��. v�φ����て�=흃�w���������J?g�н����Sa�a������ѿ,&#V�����0���f, '~}�`�8�)/�8 jV��.>���vz@:���[�{���㷭~�[ʑ
C��'@�P	�?�K?�~Hw}V��k�h�c��zy��u+����c��ϻ��U
TUhq����,��F��oo����$;|�����l����/ip�E��qh�Iݴ|�լP�����z��r����C>
"6iQ���g�q�>G{�w}��u���E����	ԣ1$4t��.ue�;P�!lU�� �F�t�<�u^�FݟU�ޕ~��\��YJϲ�M�_��;} �:d!�k�X�O���:�(
ɓ��A�<(Yf��x�/��Y���ͽ��_���P�����u쫻~\���	��͗GVל�����m-���n���A��������jam9��L�a瘐'���H���5+�{����8&ݎ��@��ϝ��K&��r����[��E��OŰ;�=\��X3���?v�M.��������0�~�հ+4y��Ed�f�'Q]o,-�߾s4 @���
�Yz�1a�� زR�-�XVV���;`�3o )�&�/�Է��㣥:�=ҧ�/O|�O�ؾ��Ea���b>������E��_��ϋ$<A�c���he�F�w�nB��98
�� cvW�%�'�������TH]�|[�\�g�.
:�r�����Df�+��8�<���Ӌ{mn�T�E�{�h��� ������<��x��)诖�ުW�M�� }(��q�?3Z��}|BpWp`����Se��fBwۘ�VU�K		��?��<	��SA�v0�N}���nZ��h���C/����[:�� &o�|�*y�o|���������v��k��_�&���P�w�P�}O�A��@?�,=��V�L��o��m���
-��ܽ��ݰ������`�N�ZX|��s!g{���Н����9%���_�KK�iAؕt%����n���tJ��9I�9%�h%����j� ,�+���f>��ф�����@��L� d��.+$��<3�4A>/�ߺ��m;���QY�FT�ڶn?�Ǘ�$����DD�?s�������KS��/�۽����Ĝ9��Ey���%���>C <,,,��#��O���8��'�ֿ�8��"���� �HuF���>�Ըu�Faq�c�r}�L�n��A�kk9�F�y+����T�ҩ��gAF�m�`C�$��Z�}�{�e{y� �X�`?�DUiSShQ�\����4ϳg�4xxx�/(��� ��o�߷��T���r�IZ7n�6Z�-E��Q_#�[m����]����t�M_όg2d�GV5�s���ǌ��4�+Փ�v_J������������洈�����:�N��d�� ���	߼���,!��ܶ���B��h9�Pp��ÿ�{�N�5�j�-�?m��\ku ��Ѩѳ�S��v6���fG��l?��M�ɻ��ܚ�U������ 
�dg��1���U�������-7���U�Tj�M�u�[���brb2�'l}��4���X�z0�����8�U�i*
�~n5e�L��NQQ
7��z��@�؂ss��7
뛛�e֩��J�'-�)��󥷶����o	�>ʮ
TN�9ٕ�v`�sKQI��n�<k���՗���oa�3��	yƅ��Yx��Pi�t����S�j�;m�#�Ù�����.�_���hj$�ߓ�����}��2>!Q4+���s)�#-����P}��OB����߀m���F�to�ȕ��)i<J�㩬�;���C�������/��mm����]����������qX��dd%K����?�����PTW'w�D��4?�V`��CS3��Ǆ����~U�|/<�c��������O�C����WQS3�np��G�k�4��"Џ�m�"3��~��
oߔl%���9(���f
N�:X�'�:ɼ�m�)#^�4y���G�%`�:9�AEE]��^�O�%l��IIIQ��4{ Z�{=��?<x'[DE���ӿ��$#*ټ�֯N����0P�]���c�����[Ӎ�/� {�ʃ��\t�grnd�r�p�y�U]�o�-0g��2F��R�ƠWg�ƿ�"<�~�ܜ�Jf2a�	U(�
ϡ�)�����PM�u�]xś2���DEQ�I��|��pܤ,���F]�x�]S��t`i�OI�x�����)�ŭi�&czP�����"y,wE����q2�є���#yʶ�Z��5��tt��ө��V9Q�׸O9��jsE��%�ћ����>o~?Ӆ�6������7_�iV�+��޾�N�R���.7p��Y9��~���� 	���ò�e����'�t��̀n�B@�~j!�4�V���@ �?%��Tڰ��%TǪ��c��PV��roB"��%�~�k�vQ�3���&�(���r�9�f�Ak��/G�N$��y={��|�w�;"�38������d�C�{ֲt��d�"�^2u-��55�D��n��L�K�s�ԁ[�����(=���[���hQ��F��ߤ� !qty�sN�+ǯ���|�<�R��ow��m-ҾB�A>�^�,۶�P�Ϯ��p�l���)tT����~���P�Mm���D!/O;v..��4�XFĚ�ģ��=����8Y8>UD���}��k.�+h^���e�9�Ɉ��]+�<i��:�%P�X3��F�"g�P������r*��6�2GX����fҤ%p<�����U�Mî����{���Q�ǋ�C�_I^���*�����!�V�i��h���kn����ds�d����,X�h���_���I��z�óU�`�\��X�9�mS� �����T;*�A����*2ى7J���ZT����@ l����/ϏW���ע%�N�`]�E��hh��Pě�������-Gd���^?�j��~v
>�6yN���Z�KRN�i7h�T����]tvvF/)Stx�W^�u�v��4���o���
u���F؟e;��{����B� WLMMm9w�.���J�̛�U44X,�?uHj�����o� �W�V��`vS�oh��Xt*Z����^�xdU���a�1;��ym�+Jy��T$ZK)��P�9`��[p�J=M�$�Ϻ�}>Ł����Y{����3=%��Ca�@y�������Z��,���MoOՏNM�T�j3�-��$!~�ў�j��hOF�d�c�<Y:��8h��p��6���m�&��B4��G�{��6t5��1:&��5���gN��w�c���k	d~u@��p��Ҷ~
Ec�]���.�99QQQ����f��!�U�/_f��d2�"[o�x p%����@��F�s*�L�#�'����4!�p�C�yu��m��e��$��n����wX�I��ן��vAi��,MEZ�C>b�Ps$38�(޳s���1̎����
��:�I��x>�b�Jy#�yϵG�h���b�P.H�u.���p�����T�[�⺍�j��Gͩ�KG���N��^��Ed�	���k�����Fv�%�Y���Ծ9 �LMT��o�6@ܤ�ك.��W,��0+v���Q~N���1��/�&F{]�o����p��&����G��s�	�'���:6�ݎ�<���ۡ��#�
PJ��$4:���A�p���z~Pf�)��c���f#��&��/��>)�`�=�|���)��r����u{��PY�j6V���1N�Bg����|��]���ڭ
�������I�z��ı�8�ס����D���ͼ˞�z��������^FO�I��pbB
Vt=��&���H�_ϋ���􈃟���̵`A�HSSS.	k����<���9I���==�	C�R�{���DYR�~��3����-���xH���Ϗ��@Hٝ��V��(-�N�O1�<�$.��&�sMM>3K���z��X����.f�+�b��N��<6�o�ҝ�Bw^@7�A�i�e�U�L�������{���+tbד�����S��4uX��C�A�\n�AUTW2̢||dr2�Œ���FL�N����w�J�c�<�",�����Q��o	��C~f��g�xA+�Z�3I�lb�Ka̰:5�1���8qC%X��絍���cR�ۄd�?)v�n,��,^��,i9���o"Oe4K�Y�a�QTEE0��6 ""RQV#�����Dz�g��$�|UUUt?�Opʀʟ�ϾQ��%�P�^z'm�i��^�zt���G��i׿�7_Psf-.~�l}��4��2�G�g{�Kc���h���/�k+� ~;FE��S��ϡ鵍�њ])�nk�Z�3�?�a/��� ?��r��A�+ �!�556��+'g��T��-~���s:)++�����%�;���1�]�#�u�zrkd���Z���_&����Y"zAɓ��0q�m��E�v���P9z���t����z~�3��Sn�v�E��`��t?�R�S�9�\�PK&�%%��I������$���=��嘘<J�Q(�z�$�<k��rHN�h����
�������*��i�-�%�c7�^^ƀ�ë��� U���hm/peI=��
''�Tn���9y'�,�a&�0�AU=�b�����zw���|���\�t��7�Z���"Ǹ�^d��u>���?���p��9󃠤�ht}���ŭ� 2P�T�B�aP1:�S"@۠n���5/릅rD#^Sa�����J��ċ����tGC����ń%�Zg7!���m������2M�F�"S�z��:5��7��ǽm�NiF#����m&e�F-o-��qu}�Wx���M_vrHH�1�y bҭٞB=�����b��.ڌ�cړt3_+�}N�hEhY�h�$�W*��g��:|��k���^j�8��c���0�/��'p��M��C3�!S�+��J�#�(�zkG1�Q�xB��Hm�E�khIO�c�-�R���լf���m�\����>��s=]��'����`��U;U����ή?�~i���(L7���|1 ;�^/��E�g�p�O��8o꨺�X(Y����*�� P�?�z���E�V�҂��L����>u��։(����%%+#c���!����os��KaG$
;����u�M�����ɒ�@*S��c�˘�i��^��mtW���8�~Kq=*)�$r�$q���F�,�<Qm��O�D����O� ��0Κ{P7e9:2b�~��S�h/�¾a<�4�(��U�fRƙ|OA�cS7r��+Xu��R>��B1�4~h(㏊�yyRrF���0~RX��c�L�(<D����ol��6�½۱��&U����G�����:�	i�P�n`�����W��Z�0w�ɕ�R0������ԋ��vӁI�)Uf$��x����L�d��h�=��	��ѥ��K�����k|B�n���Im���+�H�9ئ1p�o~P�rG����F����B#�\0Kv@��f|(��Uǵ�H:!��{��2���ɪ�|�SA����}�2r��-��i�B�_
e��T<%t.R#�_��%Y�I��u��PZ�%�� ����=��t�?�n�j��s!��J��Ǭa�j0|@����<�=�3ك���r���ɩ��a���<P��q��-+�[;����h����
��t�����j���^"�PR�d���diZ���O^��L�z�^NXޞ�5>>Um��M�b&�U/�gB�v�׈������u�p��X����<�X�4IrW�bb���J����T75	f��x����53�B��h�c+�N{���cC���-��ص�\&_�9²Z3N�1��~��A�N�ӧO./4��9���cc9��v3߅�J�o�N7���re�|�t�u7�um����8��:z��[K�<wI���e���K��rD��fv�Y�03�:�b��SP���'���u�iG��= �G�~A���8Ƿj�CuTU��'���m�N&ܟX��Z9v�с$):3��d�s�6��$I#?�?��]�>���ߨL�Wײ�S+|�n�۵D;3<e	�8=���GDBͫ�nE*�c"w~f���lT���}]��D��4G���+�uf�6��:�������.d�����j[���;������c>���,.fAe$Ń�����6ϔ(�ʥx<�?vs������,	 6 �R�g��B�?�J��m;J�j����ōG��FUm��]dx�8��W������f
�V��P�w��u�b�qGP�7�=<�+T��H��ίG�'FB�b�ފ�ۚ�M��f(!Ǳ�?��쥤��U[�^h(V_�G�G% �?9y~II5o�>�J&W�<[�ccc���ܙIN���nz}��n������/៊���(��,%.�%�P�}�P[{�f�A��_����RRW�մ������4�x����p��~}���Ծ�Nz�[��e���=$or�Z��N&'[�Xh6�L�!��D.sd 
.�&��*�)ccE�����F��~4�e,}�x�\�20�t��B�f�<'���G�>{�5�ړ=h(N8B�ɸ��'᨞��V'�!�[�����R�Jt���/�r2�+�����&�<�)��D��|0]4 gjT�ֶ$�����Y�0_]�3��$��$�?��Т���- ��@}�F�u-�-vF��ʚ�n*݋o6��U�O��p��%Ѫ�Z92�{��'��-�^?�Ǎ0}64Ð��˜���2\�;�?p���"�-�&&&,���J�װ�]p���J���>���A�Z���S1��R��Me�館4������ 5�#ZK�߳�{��� O����t3Z���`����ju�8�����q`�;�.+�Nr9`�����r�0"]��!��y:mҒ���BA}�q(�̿h�D���~�}=��Uo������E�Lj�K0�2�{0'�1
�G6�e�a�b��n%�^W.��=HLNN޿��w���y.��\��-%ؙ���:c2T�4�~���`����u���(-gy��Hz8��r}��(^$��c�d�l|����oky�VW8/�o���~JA��^�\> Y�
֒��v�ڑC{_�5�rٿJެ�e���&�u�V9n�����v�ceu5�c�%e�����ˣ	�y��A/P��Ō�#?��hN��G�;sGm���� !�}S����������saBN��<d�Q���{�o�A`j�~��h���B@@`}s�w<R�(NR��w�����xy�9�M��#hj2W�����{�{���?��) ��~����a?-ud5x�o��3Ivǹ���K��5fe�0��)Ǥ�B��A�	l�Cm]��f��oB����S�Ǹ������g+P9uo����ļmq�=5���޲㌣?J�>�%%�P��d�3`m�&�S��5{�����V��"A�vU*jk?���J"NEB�~12hu`DTY=���F��CRN��eC�&�$Y�S���mm�����=X8��<�0�3W���X�
>_�ݳ�s[,�w
��@0������ث�e��v}(r> ӳݎ�� ����F��2�r����P�����&SC�}y3jy4�h�~f�'>ઈ��ENC~�TF�2�r�]�����ӽt
�C��p2n�Z����@�ä��$���UϷ]#�{6��Z-�p��+��KX6�	�	�p୭H-�_Y�f�:��a�J�d������?磀'���D�����T	#�������8-�J�:m��:N׶���܁����W�U�i�e��E���:M����?���*���!��V�I=���VvSSh+�Ϯ��	0�H�S���{���9���SQ]�e)z�0��5���lg�ˉ���	2��6Mu怭6�E2��4��c�BJ^�~�a��f�Roj�aKޠ��*��/���M������,��x!����9�{~�� ���p\�WݬJ�Z�x�f����É�LQ��kd�3�71�����K�l�N��P�BhGF��X�\ҋ�~'б��2��EB��_r|E�Y�W��#�0�����^Aq]~��5�d�hǧGT)��m��������s&1lx���<�d6ڐi��h�t[��C6 ����	k�|4,c����+	7'��x47j-�y
n���8�"t�%��0���
,���Z�L�X��vz��u(���\���q���g{ˀQ�*=����������^2��5������sv�k�ܶ�]��ܯ����зڷ�;���&����!���ʑ����Gl����ʰ�k�\B�%��y��+�jj�P�R�rM�l{8ƣ��5��~����]��|���v~�n9�k`T�����`�}���*�O%q�(�.�z���ߟ�O�1�e�u?�
�ݩ���� \��b����`3�l^圈؈�%�W�t�_?�d�>�w��������h��s�-�ɼ����	�P���s�ig
�=��ˤ�(��S�'���l�Ar��7r^�l7����ѽEù�	Y�;ѿ��BP��HND?�n�y�ɮa���X,����Ƴ�	b�VvY��ᢹ`\U���o��'�k*'_�ɗ���H4�9y�wY��r���K�u��Db�zX������ݻ�h����&������[��:Y�e�D`_�b��M�K�0����_ǋ��L�
HH�w����"��:osLY��/쏞$#܈HJ��3�<�z(T�5DL��Ie[x�v�&�x2�8���s��J���yyP��z � S-}�I��EI�U�e���{[�:+�׆��V��W���&��,Yw*W�ṠJÓG?�h#�ĕ��A�r�&\�d�dڪ������ o6K��~6���K+�$�P�[��W���<1����X �K�o�w��*���*v�����8�S�(ZJ��Cq8��o��~!}��H����-�Fhn��֣1E��G̓OdP.[��Ժ������������}N����ꂪ*��q�Յ 	%��rF%�`]t��蔡�ў��J �?+EQH�%w�L�q�'�)�9�%M�Q��d]B�8�:�9l�uY�:���o9iV�a�3�T7!>��&G���g�j���(�9`k�?@��%)o_���=�NV��s�o�|K }�,�`C����lc���x@�C�h<׿�˅M"�l�z�2ɹ������)K�u�76~�҈�kT`A[��&��[[}�ǡ��>^O��'(�eߣC�eX1��w�7ӣ?%IRyw�?��%��sQ7�Q$�ht�Ӵ<>����#�����]��p�n>�����"��vގ�n�ԍ?<-�����̫���":D��F�4�����J@T�$�)����"i���%�L���$O/���ᛤ	ֲ���._��n����Q�%ȷ�����]�~��b����_��ղ�e-I��t��,��~�9�W,u.�{�9'�\O��>̷I��?��ke��}u���_j<H�qT�6
��>�C����^'萴K�a��0O�Ϋmń<�9�H
�4�zU�ʶ�J�����H�y41������)/���6���o�N]/��h�8�B��9^}m�a_2x�F��N�
)w�pdQQQ���������
�\Ff2~>n&v�I��a�C�=[u�7�3��Qo/�	��]��?|�-�cX>n�U�1�c wL�TXc^c����X5V [?��	����\�,VɌO4ҫ��h:���3��C��
&�F_6�����O��0(�g���H�ݮo����ڴNz�<֯WbCJsr�}���/�����@���+{��n�.�:(�	�M�~#QQ�9����ϧ�$��V����x�g�E�^[��M�<)r�?(�wZ0{�s`�G�PcyW��	`����.n+2��C���$i�w�r�D��7���3���#6v�<,%�z%bz�ֹz>�ny	�%OM�1ߵ���J��X�᷑��y�d���i7J�J"�8r�(A�e%z�� �t�t��c��dq!&�BͅQ3��������Q���YIcU��|�H����e�Rc�ӗ�'n;*�/�G��Γa��k��-�:VV�/]����)�$���������j�c(�j{�z�g[?�_XX�������I�ˍ����,\^6�I��{]�U����h�d�3�%A���U+����c.���k�%�����^#�̗L��]
X:%P/�u�G�?\�ݵn{]K���s�c��{̲φ�E���.�����;X(�Z:D�=��3��I�L�r��]ԥ��Pߛh��ҔV.y��q�:���ڭt[
i?�
�W~v�; n��)ϫj�%�ĉ���I���$/�5�'������n����m�F{��POBuu�Yk|� Ql������W��Q���i����t�c�H�F�J��;��$K�!�"�EJ��妛[ x�ё#X�Xg�b����Ԕ��qx_��V�"������K�SҰ���F$=j�qY�NfQ����� ��8-��;��[0�-�l��,�R��̲L�@��>j�R���c?*mQ���#p�߯AϞ0��H\Y�k���_4=0�@t
�z�M�px��^y:Qux'�La���{�8Tj#�\D9B�耹�98�l��q([	�~������c
��FEk�~�Bc�^9���>��i�,� u�}�����A��ô�Z�q�{
9@�fB�+�b�-{��n��`2�?�K��S^����H�9�	��`�]@$�p��p�T��t[�$�Q2[�٩�`�B��
m�#�t}�<��/��o�5�X����a�s)?�i�
����g���2{�i��zT?���08����d��y-�ԋG���@.���u��,sG�a�G�������V���:~�1������X����e`��<��	���@3��R�յr �y/��y�XHb"QeE��� �0�rG�$�ϭv���Y�|`������TfNw�r'����,��G��Ρ���MW2Rr�����G�u��l_����j1���e�Z��T]����t>z^T�0Tqh^T[�3))	#Y�H:w�W�A���Lɯ_���E�������#^�X������ⲥ��Cs��7�`����$�/q���غ+���Y�qε�J�,ĺ��q0;N��y���`�� �}��S/�`�K��U)��+�i�׭��l�9��5EO�d����W�<�{�zu��n'���A�Ļ��]�I>���>�ʵ��"w���B��b�o	ah)�YAhKM�H�PV��u"����"2rl�vC��X�w	��/���qh(��ȓO!!8���sAt�za9V�I�!�i��6����Nua=۩gy�~������'�ڞ1�,��X���1$���!��uo6Ԛ�b֭E��y��҆Vل�at(���朣Sj�;ZFE�{M��.%�H�<i��{�S��<R�ؔM��]q��\�E�\ta�_B�/�\�-O:�F�-\^��kYzU�[lI� �7|-�iZ����RdT�4j����	ͯzyU��J^)� L#+SSZ�����\I�Ѡ�^���ia�/9'+k��?*��xsr�9_��H.��x6/� C�g	9߇�Hc�8i�� F&3�}\˳��2���t��ȋX���l�d�I��e��ȝ�-����PH>;�nf8`�M��M�eΜ|���?��`8^۴�Q�Ӕ�CH� ���p��I�����v�����E���eSy��us'�	lfp�ɣ����y2G��J���_�����6�FF�
v��Sሂb� ���am�4�V�Ы��C#��^,��D2�]�A�<,��&��x:Τ_^�a�k��]�4����\�2���ܴ�Y��?��o8:��04�������*?|^�Ѻ��:e�,�,���r ���T_@D!��,@�G%����]6AB�3`c�ZO-�#08��,:�#������c�T�.����Z<���s��kC����֥PCi U��-�^�;�B��b�����e�ٸ�'�Q����]��6[��Q��,ź����6d�W�3F�T]���]���ְ��̏��6*N�fT��5H�
~�Y�[��W�L�\��
"&�b&`�v���^^�o4���(��߿�u��907�����W�(������
�ngg��6�c߿pL+�NN��-;�6K�J.b�eK�>'��G߮���o�u��[��^���6�=+�������<�^|)���j?�N��9D��a��-��������zi�1xy�d�Gɱ��Q��lV��ٖ����ؚ�~y�z�P�9����Pd���Cd�k��W��l��T�K�8�x�m�&�9�p���A;��*^��,��ҲX�$���>Ȅz8�0�ٖ2-e��RA�A��]+c�5ȥ����$y�L�iK���(X3��L�(>�`�h����~���)y��EEE�Ke�*i���+"22��v2�ttV�2�q<Uw�k�U��X9�{W��C���5�$���Jt��s�c��梯;4�c�.�����仜w��J��~[o�2�Rf�~|i���u�{�4�-���U��q�w�{֟��h��(4B�T��0TA��^)�k0�};��]��3���y��C,��m�삂�t%J\��m|���Rmm�֏�]�fݪ4��پ�(T���5���YR���ln7/_�s��y:
��*&X�\��j&�HF!��+�؜�r��`(���ϩ:\��ٝS��C%�y.+.�U�m����.��Q��A�/C�c���D���ySc7�s{�KW���!����ŏ!�ێ��N]{O��t p��zF�B�H>��3�׾a���m���;a'f�yď��X���1G�r�ix(Ǒb�$�����Fm'�S�U�\���&��WWÇ�z]'�~��Bk��|�)���p8���c�A��;��y����������ߟ���:7ȱ=x��wc��;J�0��q6/��QX�f�.���U�L�y^�7+$e;2��G�[@Eټq�4H� ���tw(H7H�K�tHwK�"�t�"�"���]�����Ι{8gٝ�����uϘɶ�E���\{�}�7�4Y���o�o�;�9��]���Gy� �B��ɭ�i�� p:	�G��Ղ��L	]�csu����MM�"�����\��^�Wb0���Ƨ)�Z�P��|g��x��o�F�9�,V�ڑ�����{��ԯ|��S<��orF{����A�+��^���SMM��S:B��)��px�M�*X���Z�TdR�����I8�kR�rL$�'j:��U+K��e�d|�}{��2,i��÷o�*�5�x򦿫6y���:\��uQ%��=��OÆ�5��]O]�����T++�U������]������UW��zZ��B ��ϗ����"c����Zb��ML�0��⣣�_��LxR�O���в�7e)�����r;$�Ǌ&�����i�2=+>֞:9;������#Z���  \�d��'�n�����u+�����N����G)����������z�����P�u{�<e�9�Q���NMܼn�R��m+M��M��a���"n�z��x��Fa��F,ӂ�����D��M���#�Oƪ�E>�F9����4�j��Q&�u�Tk&�ͫئ����T�N���Vk=Ѱ_RR�jP³L<L�ə�"={�E �K�{�"0a�=���n�5`�LMԎ}����2=�~��@F���x ��\ӵ׵�w��ATE��� �%�Fֈ{�B)�?W*;���K�V���/�6��M����SN.ZԿ(t֦�L��]�E8s�[�iH����]b{�kH2:
�m$��I�foZUJ�h�Ij���G3����K��M5�Q��yٲ� �Ju��e4[���",#J�x���vc1{@�6�ʜܲ� �;���-��{f�-R¥�[/�L�]d����|���[�:����02�Ҥ߼W�r~��[����U f�
1z����F_�֫!�=J�-=!G��u����Ϻ&�	ϯ���TÉ��'��!OW[���}p�A� ��	䲠�M����c\B��ť�����a��z�7�3�[qC�/�D��R(�x�:�$s����tx�Ջ}�(d�B��d���q���8���ʭe�������u�v]]lS�m&7<���W@I5ߟ��W�'��Σz(z<eR-�|����)��\�<��������������ޮ(o���[�)u���cqy{�����=t���l��9$0����5��WR��3G~S���Ho�{�LpK�b��Ȩ:z�~9cE����*���ɿU��Ըc�Z����7SJs�_�GӢ6��n,�O��!�N#�ɘ�.�!�e��?[4$���9;]����M!x��~��X�Os��`�5F>�Kz��'�e�^Ђ�Tc����x���Oy���mf�S�2��ܟԒ�����3�4@�Gɱ[�$f���ϒ��ۂ
��"��[-\	���\�~Ϯx�R][����o_�� +r���1��_���*;��la����{Gr#[�Q"�����vѥ��h6�����#|w���"'ǲW��,������ �Xd�V&&�kڟ>�e*�V��������K��J��XM�yg�ۨ|������B�Q����Յ����~WW�f�x��/R�gL�lYF�X���'�'E�p=�*�W>c���fs�{�&#?��$Q��N�Z~嫝���N����k�֐︕z����T�8LhV˲a��]�_
k%�vB�Uz��
:���,p+7J|sx��t�� �ַ�1/�sǽP���sU��������[��O�j��_I���]a��=Le}�gN�?L�T+RCdrg�y�������_��Ԓ�H����VT(�
�E�ک���lq� 	1���ַ���w]t�V�!E���p���8d�~���������Q�:�<�l�����enn���"U���z�!:&f��[Hy9��V�X���d��(((t@��c�~�����p7��a%��Z�MS8ꦭ���z��H���:4�imS���W�o@��0�}�qwuq�N��O��	*���i�
X��+a�	�1C�.f�3�,����?��ba��L�]��T�z^�Z�����"*� p�{j*��@��T�5><�Z�0��q�( �
��^�}�����w��4��-n[������xDRo�\���|��*S��L� �9<��e�X��s֢Y#G2�]"�R����f�k�z��ב6�Z�Q^P��I����װg<c(E<��f� ���]�����f�8�k{�B5��>�j_��vfQ�@u �,L�a�'Kv/R���p���q�HYۮ���ͥ0����7�ګ���LݎV|�{�;T*99�x
���i>�!s��H%�~(��iJ�/<k�V�e����MX��.r9���G����֮D�_��͵��+m���A��&��k7�M�벏�B�� �ʣȷ��DO�{�U��	n�׎�ɝ�l�ií5��,~|Vũp���ם$�����������[WL���_k���L͵[��O[l5�2�Gs܊�����S*@\v��ŴQ�D��Q9��,]ڈ�F�����xȥ���K�l�Ҩ�����G8�1:?~`o�w2<�?�{��W���N�ͶKۑ��N�Q�1��7�3't��^S0�Y�
��[��-��ބ����"��f����i�QJa>�h��P���I����v1gљťҵ�G��1�����?<E���$x��}N�-dn��'Уۻ煌�m�~��?����΀��u�~�������l�h���K,��`X}.&!E}Gd|�Z22���O�>w��#�Sg�Oj��l�Tppu\/��^���\�q|�z�^�$j��sI�O8��ށ�Nv�tb�<�O+�u�6�+�.���>���?�lM�\vJT0���Kl��mg<%yS�TaV���w���@���ˁ�ҵpip�; �?owkhY�bf��kh���N�Rl`)Y�i*����eo~^���GŌ� ��E^,�UU-�Ga�ށH��%��t�b#���U�����{#Y+I>�֤]ta%�T���9�tr#���3e�D���Z~C`3X^ET����a��F�:���� ���zd7<����6���ԛa*m��k�|�Uz�Ӽӂ�|!�A������YvwZ$�uw��L�C��yC�ի���k2���=��i��m�͙t��3��;K7#�N:[,MC\�؇\�d�j��/Hd�>.T��^���f��Ȩb``���������0`�c���@`=�>^V��y>�-�\0�-�)ɲ�I0��9��$-$��ejxz�_�����w;�c1aG:l�zT�?�����-?����S�S�xΩ�Kn�(����y}�¼�:��{�gHhf���:&�
|J�釣,�FN���CL�ﶆƇ��*R��nw�۪���r��]�BԊ1�2���A��?�*uO_��L�_�2���a��lU�ҟݒ;���k��u~�ʪ��a��ɗO�Ƌ��(Q("��_��n�H�P���lL0���,rA@�8�2�P�7ӰcN�RM&
k���.w��Jc5b �Յi0�K��v�e��0y��"z�ud�8͇��>�]e8��T���=�;obf�$�R7x����c;EMd�C�q�T�v�Hz�,��X���p�ZׂR�����)C�n����բ�֬3�j���Y�w��^���T�l���'w�t�����ǵ쯇j(e~{��im��+���@h��/3T�IIH��z�"N��U�9'�KS7Q�Z8�<�^�
�յٳG�|Zy�f�4��z���!�s�`�w=b;E�-���?�8J���������kz�д��[��A������piH}�t�3~������	��5>O�^u:O��]�Fx���U��$b�,3YJ�,�_��[:�ߣ��ݮ���R�k�A
�ܭ�eCp^8	}N�������MMX�Iz?a<	mK����+�-�t�r�%I$P��2q��ڡ^af��$1��L9$�K�N�5 �9U�VeU�m��O<�����o��a�
P9ac��{�~`"U�R署��0!h~qR"��#�~����V�.S�\�r����b����O��%1�@�oUUx���"W��U �,��=GG	j��yk�qMމQ��9E��k$3--�?��{	�E�h���i��$G���� =Y�)sp�}�H�����x�]���K9���q$�߽�����GO��M��JkR~b�}���i���t� �V��̘%���?��6$>�D��6�������j�� r؟y�� 2�#�*"P�9���G��v+��B��؇Ł OU��(����N���c�Z��*����P,�="_>>�f�;�8^K�?���]&2���0���NQZDo�z�N}4z|���;��$�j]�S��~Z�MO~o�j��q=�Š%e�.v�X���0��~������,#�.i�/�*]rK�Y�Zy�G��}=��cf�7�o���А��4*<�c�1^�d� ��wq�k�����+ה�qg�Z^�YQZc
p�'�d�
�hQ����ػ mˆ@fj,qΙ�7/<i��-E9G�:�c�?�)��÷�a:ޘN�١�\��g���=h��f�قV
�>ڃx�h;|n�S+XlA�M�qT�M�����ݑ��W���i��18p�Ә���͘j�[z���e�?�|�cy��j��Q�uj����WF����ă�@�,0���&���S1-�Ϻ��{���a�O�����!�h9ҿ�Z)��ـ'*�����4dv���k���h	��x�e�Ǚv�n��n=2&������A��f-���~[�\���d����?�[�߄�#fe�R�������-h;Ƚ�o��/A���"��~p'L �fL��&�H���@����gv�*����CP��/ם��>/8tam�7gZs��	猦ډg2}�R�@����/����p��(1lj���}�Դ�F�Wh�M�P?�Xy296j�!;6�h�A����U�n�Ջc�FG����|�wf����5Ͷ�ca��n�>.҄^������7�6���Է��Än���j��]�FM�6�X�:Ժ�s�A�Q#zBBC��
�`Q��D�jX��[8�kM*++� ������P ���W�lZNEOxB���(�Q	��;�t7�sR�2k.�Ӯ폂܊\�35�A�[]i\���5�~ch�J�h��̠��D;GqѨ��A�N�Nw�c�zSPh��d]�t��O�Oǹ+VX�m�>�����a�铻/
��؄�?��B�H�3^5s���q+,zW�a.cڤ�]�>�Ƙ�n�鹈�H��tQ�O�7Ci\�|�.�IIIK�zqey鳙V���ҸHh&��V��@"���愤�������N<��5���ɒ�'�o��f�@CB &&���I� _�;�Ķ�嬤�X�2vG�/���E���3y��.[ޗ��/�ڒ���,:�S����`>\�,e�~��aa�l�X�~%��Ĳ�H���ܮ�=��vz�N�VVV������K�g�ܼ��>D N-δ/]�)�zcK�z|5�$�G-jdL�����H�e_���E��#|h:<��O�:��Z&����j[��[��8^����E����,�Ê��[Ea8lW����k1�X��h�󛶥�M^�[���#��:�g�Z/����7���޴�Tk>-��������T�>�r���}�%�_�\�Ч��r�LI�_=>>ZS��������c���28�g�Ib�Ј�Z����\�����,�����v6o��L��bF�d�Fv����j̜�k"O���z��q���Y��@"#o<����C��yy��{{M���KQ��^���{	3��m^�f6�$�u�*O�ﾚ�(���o�g�T��M@�s� �E�������8g`�݊_tz��R7���J��OJ�+���a�9�������U�&��ƭo�h"�Hj\�94���"�هP�X�#��^TTG���:;]Q\�������$��J-i�W���݋P*��{p =`�T���gu�������~t��:�7��Gz<�NB���cY�.����w�rvWlEֶ��Tf�lw���J����~+-!e�sVl\�FĔ��M��z�Lm%]����^�YLU�%�e�e)@!!�.�lV���9�]`��+���y�y�j��_��=j�뽠���e���xx�E��|�y��x�������j�K�����$�,���"���O�v(k2���ۈӈt����<|�r�� ƺ��B�2��G~,��|�v4���$�0oߎ%��)�!{��_%@G�w��(p)�5�H>�����O�~��U�����:ɿ����؃�8�bw��R��]�=Q@�N�?��S�J{_�%,�{�yOƫ$ؐkK"\R.y��R�x�6O��>�.t�H%�5d�ϡQ=�ss��%�><iu�}����YJ�����`��r�y��O�tJ$�v�r��8�,���6�WȠ��w[�6�7��6������#:�`q]`�ND3��e SWͶM/�W�h"x�U��$ �n0]�����������+g7��/J���j�"��>0��pĽx��ɋ�`���0K\\ ��Hj�����'4����|�g��ʚ~rlaJrQob�		)eOA[��xvd͐^������6�6�O^k_$Z���-jv�ʹ%�4lĴ`�5�{���?��tMeEK�PD>=f����c�<��2` ��8c�r��'�.'���#g)�����Y����F)ܱ�&t^��]��0څ�)	��b34}����.����gb����`�P�/��D�����7n����P�@I����Ns���e�؇u��W��\cI�~3d/�����Z-D���@�¼X��T�#��#YB��?�Kh��.p����nE�f�M�"R~�-��P�Yt�)*�[G��:�R~�	-���[#A~u����̜�6�:�����T~�$);w��p춠��X�˪�I�TK�9������g�qW)�{�K^�%QϮzc�)����w�Oʘ�$	���	�q��桡ܸ��^DˎON+f�v��޿K0��*V?	��ڞ�.:�2����:Rs�:,�,����B�3P�]iiSS��n�ᦽ1�J%��u�z:��N��퍕��R�?L�=�_D�+��a��~�zS����KR1{:���[ڴJ�y�9���BD�pp��%^ԑ���Ͷ�����!7��l�x�t7A������?��ц_��L���(���%��-����������lU;:����7�BJM����hU��޵cOh# \ �|Ê��w��'��Q��Nҁ�KYB�i��a�^���fl_�����^BCC*VG���� ?��E��T����B9�M��]��~J�������{�n�bu��f#����Z��o��|�t��$x��왽=�m9>U'�Ѿ^�j��4-�U�����^����nl��<�U��rd���.�}V�Wy���&9k���K�+K����Q��&�'�����gK�?n�q����@$x�a�g��?h�������qI7+B�J*�Gk��>�E��<Z���F���.B7�$�9p[�X�v�	?��^�Q�򥣴n��G\��Y��;T�6Cć	�kS�Vچt�A���L�K���G� �kC=y�Ҕ�&�#^��KI!��9o<髠�Ɍ}4�]��7n62�Y��~��2S���n�y./|� �1`ط"&܍b~�7�i��D���c���%�����e�غ8?/�9����<S�t�R�j!e��'�#�
ITS�L݉��Z^�I�S�'�7��Ȼ��"I��5�
�ف��E'j���u��c�	c�t�����&�ol�� �@N#c��LB\3T��|����D�����A�(�7l�x1�յ�2�f��Nh���ZP�^�5�U-�ʞ����y�k�*;B���NGS�
�Ю1W��h}6�i�i�ơ��6t@X�>�Up`e;Uک��	�F�N�[1l�O��O�l�{b��;�tB荈�gr���}?��Ղ�K��):k��4��E����O��b�",�s�)<Ї��^!d���=�Y�P�c�v�)E�.�q�Q�>�]�������jJ?0�3�+I�Z˽�I-Y���ngx�@���g�"��dW�Q��5(n���A�o�d��(C��_/�Og�dg"#�Ƅ4��<�i<�ͥ��j�Z��	�Hq[�ϊƻ�]!D&���d'9�����e{�مմS<�e���<i���ߠs������D߼��_8�>w�49�����gU�-�L+���F����<I�Tǧ��@�y������Y�A��,�~�^����M�vf~n����z��-�w|C�˽M
yG�ߍW�`���8��C��gf~kߝ�ZeA@����
+PV!��O�q�_��ު>�u��X���g:�����y]ϚB��D���-.t;g"�-���!bf��m:N�B�j�mצ���L���Y���5]�n�'�8ł
�g��f�gp>>>ڵV���ŏ?�kL��y ��G<���cD��Di�s��*�Ol�ZԯO�,)Ը6Q�U{W*	���)��`��*;�s0��W.<���aV-((p��ۻ��7_#[/q9�Y3�YH�SaJc����Y�怨X:��)i�
�Ɔ��>�pL��ts=��sJ��gCv���j"��({ݻ�~h��{�}iHqsy�>������nV��~��+��{T�a_̆�x�JӮf�_���,�}!�)�R�h�7H��V�6�7#�<PX�kC.d���[JV"i�*�~�☥-d�R�oޠ�X���(�u�,[� Mb�JH�ݽarcH^Q�G�7y�S��;�Ʉ���g>�$��r�)�+�|"�1�3e����(?��Y�{�??�I��[��F�r4�; u`���A�0p�F�&�fJ�l�6 �g���u��~�mO{�Qa�S��D�~���]t�cZ��c���I<�w�@�nP�����+NrZc>�nP����r�=�x��I�=��j=�u�xSY�;���>�X<*� &B�p�y��.�Vр��7I��&����8��(Q}� ���v����t ��:��h��N� ���(��I�bfA#��j�'7�P���N��D�[ ���� C�y�q�Ix�Ȑ�xJnR>! �śڳ�ꌿL/�I{o�p{�в���e���0�v���Ne���1$��*��)�^w�N_�Rs7�E��>��o85:���~?T�ڿ�S"���ykDFK+u�\噖���J�O	������5��u|D��W����@W�|����~S+�V�_M��?�i���R]�;z�\�^��N�^�q�K"��r�tΧ����	��lX�їH�]�{���L��@�7��w���nݳL+��l|>�*d><,*�}ቶ`ta�����[C��I<�w	���5Xc<���<�_�%F-sm�-P����% �8��p�;yR��`�j>��Ɯ6O��8�j<�f	q�A���ay!��E�9�e����PM-1w+?I��������s�Ol�Զ�/�m���{<��P��O��	q�H����;Us^^���+M[�R�?�_ӜN��V�;��m8����f��ַ�1�ϓ���~}*|r>�O:dZY�~Hܘ>>2͟��5G^��v��#9��Ϛ������'��$�Ԙ�,JG-�m�a�~�^�����2�݃e�as4gPL�5)�bҷu�*ޢ�m�����>CF�s�ξ�
N:�qQ�n5����-��`K�b�	�r(����	�Ҕ��t���"���7�&�7~#��a֎i��*SX%���� 5]d�F�9Z��v���D�?�9����Dx%�����gw��f�R��2`�\�О�B��Iǎ���H{wtE�7l��^@�n}�S���������LK^�ʝ��)����P����䙻��8m�F!%Y�����0����eՍ�U���\�?^���F�YQR�kK���q�A�H���d@g�z��z�H�h�h:1FI3G�+X����
t�h{6�b�F�����sw{t�+Xhd�v�Ш�}�p�+��UڥV�}��z�ۂ�o1���ʥ�B�{�U�4�G��95釸](1$��w�Ì<g�]��nI����b��f���f���p�mX���F$Ϳ`Sy�����t[�p�40dM���J�E"��Wz	E������\�o�Nə�g,>Sd:y)�(���VO�b~��{��Phx㘀�T=�v%\�fُ������͝�5)<�Ir��+薴����!]CP(􅺔�+ŉ�`*{oO4	(���]�P6́F������u.8�����F9��/zȀ��g����p5�l�&����pɪ�%��4d�>lUP���,�w��<�|��Gr��b@:���\�ݑ��Q*��}��@��ޙ�m��9�;
�<����\�k��W�<���iZ+�ʦF���cLI5=ފM��N��=�<�Uo
n�K~\�H|MQ���P'��x)�؞�QyC����,�ט����w�������c���<iJk8�X�K.�[q��O����*𽈎��JU��m�,9���˻�>�byY�0�N��	-�3�����|��cV,T4�{���n���Л�خU��Վx:�8��J�n���ZmM�g��V����|�~^�2��ꯊ�����W.�A"�aq��q"43�eq����}b��zk�Ǭ�߯�����A����Wwm�#�1u�N��>�㋓�y�k�_��|�[~�-�9p��'���mA������Kt�lE����)h����S��V�Z=�^7�Ӡ!S�������TŒl_x�24f�L��\}�� .�#'�%4�dI�/8���d��@|/Xu��gl]ڽ"���Ɖ���;��p���s��R-�J����&�缾�wS�
W��e6J�������=�w����hk�?S�*�k�]�Z2�pK������-�ul8����Ƌs���{��T�t]������o��Z�긚�'�����,�i
Ps�e�.b�doN�m��SZ5�d�O�0��%�!�>��eR�dlv����mB������M�qL�ܿ�,�7</���Лp�}�N���8�\,z~t���e��yߚ�4G6^�"�[�'�ָF n���hk
9͎R�~'�����Ŷ�u��%�������)M �����d��-�\jqS����T���+R6�&Yn��1����L�l�}l�
�l������ߘ��������>�.�o��Ã�}uxx
p�v{����`;���%qKZb�����e�@�;�R鶾�>n8 P�ʻ8�����D��m�//I�X �* q���o']�٥x�|���B�
 �H�ɗ���X�6����e}��]�3˰'��Ӗ��ΩBE8�F�_�(�M�ce�U9��#�����7�'S��ˏ(.|l|(c.ge�e�Pl:/�4�2���xb�K&]1ݥh���{%�����Em}Ո��}3�RlZp�J|*����Cii==�͡����zG�˔�����L��a^�;i�^�8zy�OO�.-�_]�>�[��~��̽��H�@���(��U��mԠ8.���~�g��-�;g�=�W���9�]�-��:j�h�I����m� #���c?��nK�\�N��<�'l4���ID������ܒ�b[��!�1}n�ٕ\��	8��n	�>���\��lo�,��A���E������� ڧ֖�^5��9�������OQ���}á�%����c3r�x�U�In���s[Qz�w0Y}q�碴Y�����/|4��������R،�h4�=@�a�n����U,�h�ۏ�����~[j����2x�F�Tvn�M�v��D{��"����DK�AC|8YYY���?�S���?�˞)¬�f�@`���^ 1����S�mlG$����)�>�(�F�W/�>
�[V%��@����h�s!��ᇯ��'�a$G,6�Q\Xh��aśhN���"adD$Q���N��3U޾UJZ��Z�,��R`{�V�^^N�@��������;;׬��abaFcac�.y'�h5�L���c���:bu�c�Mx�����~�IC;K�r[t9�J���(`��+�S��@��i���skc��Fv���}g�~�JD�u�%���'��F����.5-Ĳ�KLCy�u3[*�'	v�x"k'd��%Q�jӠ4�j��O�q��
f_�[f��D8d�?b�3u��\1�Qn���$�r��Fy�}w�i�(���8���y��D�'�\� �\���\J|�L		�g�T��:Y[��	u�A�����斖*�Uɡ1*����&�b��Oo��]:�,�����擲���L'H���EP�"�ot�5#=�����Ԩ�׎0�0$��dQ��ȓ��<W������x\ny�8l�&�hdv+����Dc�r�e�
��L:���5:����yyd���	�b�������q�<�A	A��o�G:�W�2�d4E^�7p�ʴ�nT������٥c;/����"��]54��ꁎ�/��/h\�%�s�����?�W?0�i�U���	�0��8Գ�34~Ƚ�� $f�?����c_��V\��Ǎ��N������ �f[�L����m�6)e�����]&گ ���-u�dK�.����_,������Y�칏�-������T�f~@�K�-���c��%x�f�!�e�<+C-�6Sc�u��)U��t9�t��4����[g7����\�Uh�]ͬ]����k�^�}o�gsqw�ki!�k !;�:���ׁmԄ�P����[��7�ayUUx��O�����&�zc�|����I��ǘ[}m'ݩ��6jt���^:V�4�T� ��0�3��ݧ�u�`��\�h����.MSkA�T" 
�)26��(R��ǈpC("-*�3h����ՙ��l�iqѴ�5.2����s>˷��X�#3��@#N�%I�dJD�+���� �U �>���Y5F�A�SaZ%�h�;D���0��Z�Q�K9u?�k(���ʨ�f��P}v��Q�	k�|�6�������#Z��ؗ�^_���0�����c�F��D�u���xzT�ً����$y�"���7����vU��MNjLaOB ������W�����h�ՙ5�E3�Q
'��v��"-�K�w�ĆS��(`D�'����W`Wm �:�H�,�;�``��Zo.���,K���\�di�d���r � ~�C�nB��nF�sss�l�$�P
8T�Ȟ�,�X���Ԅ��8�K6��Ⱦ6S4����Xu n~�O��rl~rl��?�"'':i�Q��l3�\9g~��+�:XX��0(=\�`�K�q���M�� ^�1}�Z\��
fӄ�P��S�B�.��=���U�8I֒n�r�ґYBo��N��=@e&���i�{.8�Dm��抰E<bF�(���=���䁋n;�Y��-��ba�τ�b�"�h`���w��Ld��֎�F�����-z��l�R�B��I��d�
�Pd���s�ZA!����p={(!���r����ZG �L�=�/�3�7��!!(,��h�J���{�B���ʯ�¤�	�Z/�΅��&O�+g	v��(�w|j*��vJ�@~���J�&�'���FO�n��R���i=�Ȃc���<�iŶ�r��E��� �(\S�R�].���|$�\�����Z�x`>�����E�n	��~�!�d4��|Ohu󇍡&�}�?K�Yf�`ۃR�����	�z�˼ܛu�I&�K�?^~��s�Y{��hmuZ]u�d��VV���C�H�Bn�`*4���¸�D��A� )d-�=��6Q���)<�YK���$��n�YuS����))�1Wg븑��c�L�_kve#�D�Wf�i�g5�p*�˓&j��R��X;.���	߫*[7${k�ٻ4�����2=&��m މ�o'+�&&�v��v�N�u.�qs���ꇣ]�V����0���e��=��b�5���VVLG�4�DsB!���2hUR���ӈ������542_l��������1��l��7�@���R�+�����ʸHܼ��/"����lmaxP�VbӨφ$��h2 c�Ud.��!�?�~�!���78��+KK����1'}�������Ss�S�p7��k`���`)�k�J�;h�(�j�G�x�e����e�X�P�����ѯb��@8��~�0��nBX�$�f���L����O:�m��8�r�$���c*/���o�\#��m�NJ��ֲ�
�������W�·��=Ӝ��1n,DRc2��� �������5d8Ӥ�I��O�вx�	~�!�f`��*�����(��B�P����J�QJr��`#)������|U�Ю����g_Q�*���0��H^{<F ��^��5��f�D,)Np��Ԡ�a����n��W���ë�G�N�P��qݒ�S#�[a-M�J�,��Q��<�v-�O��L1��yv�TXe;��
@-���$��n�*�@���0���`OP��(�/�%��}���F{e��7Y����kҗ�4h���d�8Q�7�����R�����Gc4�υ&ma�\���o�����q���\&X���
�'iӈC��:,,������"�{z�����L�+ƿg�݇�o��L!�~Ǝw����>�4���%ڏ�	-�Iǀ+oQ�˔��#���������&�ca�4y��t���;�?�W~�����?[��u�߹����*����)����̓[�wFp�ӿ��j��=�qT�I�E���k�Y^t%�T�-
�(2���+ݚ��+�f�C���Xx���,����vx�W��Ayzo��O� �%���چ���\����#&R���"�m܁�K;W����]}�9_j>�O���i����
�to�!�:T����IZp�_ǎ߆++6,8�}�;����=�����g�n�#i�}�4�"i!d��|=R���(0��'��TI-q�xؼ�0���Q�z�d.�+�|��c�H��T��!�"êj���#;���W��A^:���e��-��zΙ�	4��i�HII�-��N���8��mf�ˊ��f�xU�?�0z\!2�'�[	x/������{>}r勲6����t�r�{�EFEB�Ks�󬐨�~z� �z�Y�W�ŀ��m?1>nkkK0�J��[��;��Ǯv �Z[�&o�,1-G�5kd��ǋ�{�skn-�p�:O��f׽��m>O�2�~����N���l�=N�4^Aޫo���&	@T�qBP5��`�Oa��0�/Mv�9W���}��>�шh���>��F�!	!���������s�aBP�at̪��ls�e�O���2=�[z�7�T���q�N��Q{�� P�}n��bH$��n9M�ǔ�[L �ۻ;���������7G�/�z/��b�*�)���a݃�W�
��߼�	�O�>m��ue[�C���3���Y�����]\�m��x_0���r�ָ�5�I�,�)bK��0~]"�e�~��5��׿�Ѵf޳�ߋb� �AB����)¢a�W�|(		�]!���t��3�+7�U�!�� Y�.°����S���BjZ��(�7 ��v`Z���V�?I�w��'I��ֈ�=�/�v��K��Gb0�[4�F���t�p%N�kM=t�p̫��Z	\���A��E � >�
z�3����˴R�����&oA*�ccp�X�lw����CU�i
�\i��v��) �=�O��F��19�ϕj�\N��nM�Q��t��|���z��Z آ/�)N~`���J�{l�ɡ����畦�3s��?�|���.�A����-��4��X�Ҧ���v����3�J�a���EM���8���8I+�g��Y��^��N�C]�	���ThJp7�"�\:H��	�ѷ�WU�����w���!��(&&�d�Z��ٹ��˅(�H�܍	�Tcb�I���O
�l�aE�Q�*ue�t��_�X������:z�Zo��m����/�yB�o�I\J����!ʰJ��֒AjYD�����~	܏�`
���Uߐ�Bi�R�&|�6
�"�~׭ؠZ�[�ȧyu[�7��ء[˪� ��L7,S�)�!Lq�,hh�f<�*��.��� ��m6�p��#�D���n��Q9����H0��G��I]LZEZN��fD��8�͖���S�v#�in,�׼��c�@|��a�oĵ�.�kNjf��ΰ�v�А�����l�|^_���u�������ea/�|d_z�̮�*�chW�>���133���o����xc3l�
ņ������͘�e�Y�@��o�yf(��.W�����ʆ�m���j���/��.'p~��[�+��B��L��%�\3z�-�r~�(S���&M7E��[��|�B��?�3����,�����7G���^dN�/}c�3f��Z03���}��u�����v�q3x?��԰�Y�YY0���ͤj&J� ;�2֒�l�p
��Vvv�^vV�!f��)��.���@�<՞y�20 b7��$Z�ʹ��]r[r�[|�#���<�-F���҆�o^4n�Ko��u\��������6�&Y��D��j�J��l�ֶ|ww�֣�Az�*�?����M)<v��g�'��d�}����[D&�F>^^p]!@�o�Л��I�ߺ�� ���%�NK�;׬��E	! ܲWm���
�*����/ݍ" �)� ��"��Ҡ(H]����D��A���;/���1w�q_߻g���ٳg��5�T�g{݈�ϟ��:�Z(��jU�T���)��߂��WJA�0먉83'��'�Odv��u�~���-_V����Q��ܙ3U?�xy�[�
��k7�������!�5���f����Xy����I'E<�WW۽𶴆���G�A��1WWY9��gm�h�:t�����.�"hRFٿs�����ď�f����s�v��)gc�B~�5�eH/��p� �'œ���� z3^��
�h1';��;n=|K!�J���Z��ݧ�5����1�o�S�f��{Wҁ��	a�Q��6��p��m��HM�S]9%%��SV�c��Ʃ�#�h�����z��)�̬���X��q*.�<O�<��������
�a,�0�3�t_�[?�X_j֛��5�g�����K�k��qO44K��$��NE�П��-u�_�D!��[��$�'w��=F��;Ư�F���A�՘ ��	g�IZX�}{֕�ض�� Ha^��X1müX�z}����7s�X3�'O��0��t�^V2���T���MR�O4@�zA����i-�U2������_�9��v�z_s4���Z�^W�	a� ��,.�zJ�Ȼ�)xT��,�J#g(!� � 5��db�>@����, D9I�����O:[��.�n.j.�����*-�uRw��X��p$~��i��$�n����������t��i����	�����.�
Y{�Z~�`k������R�=#����� �ڭ��|�?�1�`����;}�d��St��̳Z$;��t��唜-�����]e:��Ч��ӓ�����[�P1��&�PE�f\Q�e~�l�H����3>�a]e�F$�|�Gq!�y���Ne��bD�j�8�l�$�hW#7:�Gm��Pބ���̵'L/t=�)��;g���>t�})�c�]��E�6"qCΫs�U��ϯ���ï�ő�Y-	�Ǐ>�),��p3����.���ֺ�/}+�!Ұp���B]��x=`	�f�e�	���B�i0��ˀU��9�6_0�v�fg����ؽ�2�VR�-�?�s���i���T��v�}�����Ϳ�B��``���D)�yA��<,_������M�Kꥎ�5�J���=��W�Ax����&�XyKA�qn�o����#��D��j��A�t�j�Yy��c����|��$i�ae�G�� �� ��� t�V~0é�1��tL�'z��H-�F��Uu���΍���~�aאˌ)�Z�+�=��w�ҡuv�qa�]�~ w�7����4�]��V��U�}�I(k�F�����}�uT� �D���=�����ā��^F�3�����8���[��E���Ʊ��tHt�O�~7
^M�!��� ����h�u!�h��P_��:nM�����v��E�W���H`xG�쩻hף�1z�����YYL��+$:X1�t�#+�!]4�g��}[h@��V�g	�h�-֏4�X��z��y��L�PU,!!��֙DPx��
 ���E�Ǻ����!�NNvwS,���?��P�X��-�ڕ~����є�� �[��qzͤ݁�����A@9M)i3�o+��.%%�K8����Bw���ȁdӂm-tJ�)��P]�ǀ��F���Y�	��_�)!G��\�a�-����9k$�zQP�I����@X�`,I�3�w�F<tz����bɨ�QS��Q�\j�ܼ��hR��n~#�p�	Ob�>Q��^��	;�S�0K�S䖎9r��X"!%�뿋��������Puk����`Dp�1�����m��F�4���,?��޻
S�w|�M�`�p�-De��b����%`�^^b`Q|[��O�3��{޹s�t��3�*��B8/����a������&�&rҪ�|M�.�{������,�GB�/���-��<�Ѫn9���5l� �gff���S-�8tj^�\�|��v�!��i�G��ܐ7a�����p�ef��L)�՗�$E�gϰ�u��mz�� '����SL1I0�M�G՟Ϭ#�����b����G^�$��uQn���fswFj�f`����lƉq\��1�Je�̸�]m�i����8�0�F(t����H�љM��1�5u��IW���#�{�fo�O����p���#��Wl���x�1T7�l{``�Ǵ��Bk��o�tf0�i.��`~  ��>h����6��*r��U}��QXXx:�"�]{�z�q�_��՞k�sa���2�����/����@�� !3�L��p{��f-+���D�Z<�]#��jr�y�驩�2/i�;LL�D;�57�/�m#�h�Sa�KHL�]֑�2w�/�� ����Z\��I�W�7ݰ�hӟ��~�*H���8�OɿA�hP_��k|����g,�N�)U�MI�ە��*ܛ96��/��B��d������%TU���W��uՅ��ST
aď�)aI4p
Y���v�߂��9Q�i�#�+6=�V�:`K�;a!�?׳ޗO��no[Ae����i�	�6����ĝ��&��������M_P�V\���n��yyy��}K����D�}�~�����P��{��^@#h�l&�������;廉�E�pݫ��`׮J-,�]�5'h1�(VI{�2�ూU��#f�3a���S}�Q�tl(mc�f���`MS"�>�~5�e=�@Ks���=����j���KQR�A�uW��4ך�R�n�{�=9$O�|soϋh}Ua�ޏlBe������99������#��4>Y���z�L�������%��)�eE����9�iшl$̒�'mW��|��̡tW���\�2�t��ns{Z^����٥��k���Oũ�{��\�Ə��L�h��r�?3Ĺc�Ԅ%/���`�F��= �4��r�x��t�H#�U�H7B;��̺=ڮY�(�=PM���L��>����Ђ^I���|�ߒ�a�3�A����ڵ@G�W���К��z�E��׵���;:K|��~i���d��E���b��ۭ���*S^}�Z0�������guRRXS'k.cc���8�z}� k�%����v(�ڍ2�d���&��m�e��P�R�vq[3�N��ԋ3�3!��8u5�É�6�4��n� z�}G�a֒��yc1_.nJ�V��C�o"�S���7f;�ӧ�\�5�4L	������A&g�~Ρ��*����Z�ٜ�Zu��+\4��b�Nc�F������ޙ�|�����R�1�3sԤ��1K�1E��+֊�����C�w.΄c,}G�9jJ��(qN�ւ`TUS[�u�i����T������[�#����0:�!(ck[�7��<cy�з�̯��N��qOO�徔��i�գ��K��$,�=	�����ә� �Gߣ�q2h��R�6�HÝ|�/�/�,�a w=���H�A���;m�|�#$K.æQB�����0��"��#�;�Շ�_~��I�h�R�|��̋>�"&Ts���'��̣@�F��\�[��a�[��冕Z����.�8͵��R	���:�6�J����frC8���P�~��Q��ɘӴ׹;L��>�b�s����feϗ袕$�����w�׼��x���Hf���ˉϷMJ%y�"'\�X2�^�B��
���{�Z	6t�A�>c�\�3W{���+r2�GnU�,##��6���f�;/QQYٲ�r^^8�6 �SSF���Z20�e�������}�L����'Q�ݙ���r�:�k���<�������-��~���JK3�ѭ����E^���GL�^���+k�$��i;��a� �Ԋ
8S��1�K~����n�%�+����[��s�-�]���d}�F?����hi����\YW7<4�I5�KLl��o�A3 �%��q_Y�P2K6��h�'Fk�l�{�dl��� &����秈�?l���mL��;�]?��2���4�J�Hܩ��A�cu�p���������I�Eo�+T�s�-���%���\}�cag�1�}$dt;*����V���)|4���˚��2�b��-޸�8$�c�b��<y�o��+��Q���B��F�k�w�m�<��T�O�>u���P��5�#''�����@�ʊ���@��p�Ǧ]�F�9Da0OGIG7�G�]�G�f���bDf���g@������5ϲ��[�4v�&?<	�Y<k��g(�u���MXF3et���W<����%�����>)|����Lã��]g�����T̰��8]�t�T��\�	%e�b�G��V��P�E�M�@ Jn�.a���w.�{�4'yS�AB������W�K�?�ؕ�R]ܾ�x��r���8HF�g����IX���g��W�N
��e^��)Q�lQr�����k��c��CS�6?ڴ���U�+B���E.je.R�M'9���^@�F1��l��`z
!��8�oLL��z8�V�qӆ��^��� ����CJJ�2���UV^�707	���+�������*���G�{����%44ځ1>ٞq�-�?>N���wQ�U��>~oX���Q���c�I��?������喝��I�QjԞ�B�0j�Ǐ`�8����K�t�ӊ�����~f�� �e������qK ����|��|r���?D��O��Th�[��b"ʔԬ���˽���y��L�d�wOr02���eB����3S�L]����Hj��˻:�����Ҍa��%���6�S�5p��X��D��ê�5�K��F욋��B�&��'g�S���J����'T�����{�Ԭ�b�)��o��
B��b{S5�2ql�gi),�Q-,���P��[Mr{������b���+yy>�ԑ��ߑ�W3cE!h������)A���eM�{�C��B�p	�A����^A��w96Y�Ⱦ87�k?�]w#4-*1]]�>�E|�JC���So~���{�^����Z= t��L��<�'���Y��ﴏϿի���(�\J����,�L�U�9������?T�K
)�C^�`M��Ϧ ;J(á����5?�r��yXo�7!d�!**T���%�'�LHv�Z�d�sՇ��Ž���3�C+OB���	4oL�����g����3��uW��̹���?Ny�z>�LO'��M~�.:xN�U�H�M�1�N��'�Z|�s�ovl��o�"�χ��$�%x-i-5#�f�'r�'�$�b��������o�����oGJRDB^��àr!`�SũV�'k��ЙŪ��3����x�4�Z�-X7���({��)�`+�`�Z���N��K��E�K��ǚ��(�*!5�e�D��xQy]m��c���䊖~<j�CG'x/|��E�����˴ՙު��!����G����5��O{����Ѵ
�>��~����%����s�.�����̃_i��jz���l�)Nc>����s_�F�NH �:4����+��P3230<�!`�!�Od(V�*W��oGݶ���(HeKJ����6ڟ�zV��&OJ���0���m��z�-.����g4���ǎ����i+�[ ���H��Қ�|(�Ց��.4V�:>.n>����5 ��H����y��l��	KYGG�0�ƻ�l��>���X|usSآf�QZ��_@@���3���p�Y�Ռ��~=��r����t�Ջpi��W)�a�N��ncsLa�"�p!���uH5�K>��z,��������C���,����M�s�����%�c:U�nB/~x��~_"Ǥ��N��h��+���ȠF���r�~�jH0$+���@q��YW,��{��*�lS�P[�K�g̊��PH�7�[�!������~7Կ��ύOB�,����*�������	4��v�JD��d���~`fF�[�Ck��r��y�$�ֵ:�����S[ɇv?��ao߽�NN���'�hUw�'�'�?;;���G�����F>�}7��hhh i��-[����	5�=�3 �F�6���>�#,,�9	���v�L��A���J�(����1g���F��:a5j��?�����(/��B�&����r!&J�
��y�wNJ<.�k������e�o�������h.U�uJ���wK�8,-8�?������	 W���MM���y��Ӭ�R�ڴ�۷o�'&\��̡ҵ�������CWLL̗zz����k.���Ձ���\	u��Ӄ#�>��M�G�{g}^�I�!������G����Ñ��S�y�z~q� ��ۑ��S��,�%���=_���1���fN]��kw!ܯCƨ޼�|v�F�-��o	���5�v/�_ݵ���V���)�ac�����5{N���a��m����v:�L{J5�Dw2|\ѧ�%�*��Ü��CThT�^ ���`��D1���U�1X�O���^U�|����f�[p�`�qd�P��xx)���T��>zU���K���h|��knβ��b ���\�ؐRT�-x�&Ku���/�ܥ��-���N��7H��I7[�h3����n�j4y6$��� ����`���m��r�ׯ��� ��S+	ߓ'�Ӱ�]'�8�<���@
�@>Q�_�A����G.����jU>Q⸥�ܠ�9^z�G��#�ѽz�
>�S�x �4�;?�������b�w{�n�U1}xN�V����	��a�K�;@�N���72��DB�8��G���d��%[��e�
�T���@�]]Ǧ�y��8 : Βn�����Ӹ`@x��GD�:'��GD@��:�����FFƚ��B{�MW8J�g��>���o0����1�]�_�᥊��c����lM`�N�
���Q����M^�w �O��"'(*++��QQ���M�Z�Գ�$?�=�z?a�I�ug;���I"?��3��r"����#Wh��G	`��y�����t=\���dddP��)^]9�y����_�9ƪyg���?K�m=����?�%�=��E��(_opV�3x��G�ϭW:�C�u<��|=��| ���z*���J>�ɛAH,�{LZ����eT�>[�����w��9�����B�°�y�t�[�4�������6E߂�YV�>r�sJߋfm�h��� �ST����B	���]NE�+�/�-%��^Wb���;0G������̌�R_�i����Xm.���j��ni?)	w;�c�����<G��pa�|N^����yI%%��+�	�,�%S[�VN�Ɛ���=�2r32��yB��Rϝ$T���f����aI�����eH$��j�:>z�]N��Bֶ%-OCغðУ�]��g]D��1}BBN5����}\|<�w�GiلeHJVV<	]��w� ~�VU����;��zs���|���,�<��Qutա��R�K�D���%�j/z��=��W/6�AE�oM�w�	b9 ��O'	)�4b����$��F�j�/�R3R�O��ÖԞ�f��v=w����\�M�uc�8��H��LHϴt4�/Rbo�쬞�DZ��N�O9��_(��$�t����N�5y�Gc+���e�'���҉�ЂBN��$)�p�\���`�x��m]Z,hck�=M*���m�a���3*%O~��1A���t����P,|�Y8��PF[�dYi��-�»�w �K|�g!�+3�A�%g8(D�FqS�8M��Z4������||�Ư怣�R�RTn�� o�5����MM}���X�y_�֟��^�-�H�锁�x?o'ۭU��������߿�Vd ק��ze��� Rκn�����>�U��[aҤ y�/�Qe���Ҩu焎�P��ǹ��L4�ė�'jpF�މ��x�M��q��h��tu�/v��s0w�� N��EP|=��S��SY���C��Q�-��||�E*���j��a��0��Hˍ6K�PIE�RRZ�G
P �972_&��ѡ!��9O�<��3w�$�/6ˡ���O�i"���������d��Lq#�\9��b(s ��+�� 3#���X:��7yrtl:@d*�72��P%>Y�s�c��!�n|�̸����4_#5��4�U�+��=Y��.M�g$�]Ao�4�&��_��0!�ƦC䚢�>.x���>P���9��D����Ϥa�;����ϳ����O=A*Ey�E�6��Q@JrtHߗ����4C®��Xg�W����}�m�w�5̫� /+�7d�0����KE~��_�wL���	 9JO/g?�����sW~
\�7o���[�����cs2��(�$�p~��K�?^.�ZקK%� �� X�2��
��S�z#
�ѓ3�����	��v��GO�M��Ձ���S�˛C�եS
}�97&���J�{5nR���W��W=��hW�bs�Omv.)WR��v��w���A�V����B\\6ߐOV���*���e���>��&h�;�����S�s6�i�вN��L!]S��@hj���'#W�Ѐ�r��q�?6�B�'���RF�ݠ&�e�ѭ���Ӕ���=���U��v�ٍ��qq ����ޡ��&��/���F{=,;�[[%�]V�N/W��R����]��7�g��TS�v��;s�c�TΚ���n��P8`yM^7�8'�������W'sr�h��J�?H�4a��eU��Ed0�(k�ZW0PQ��jDի�*�
s��:��-�9��2��5��}l�f�@�huk+i�I��u|��J��I��xER���T�JI�̎�F	1ƕZ���r�ʴ�ܡĮUi����G ���#i{V���>Fď�_��1�{���m�8]]�Uh���s�֛!&�����:��89���YB�~����x�ص@\��N�		h�NkQʘ����� |����8���OU�`��M���W�k�k��.� ,�U����ee1Y~ol�*��7���6��FKZ�P����բ0֏t��O�g�pT�����(�ƀ��.�	�ĪP+�)E��U<[��9��m��<�k���kg�1�q�vS^I�r-���3��DSP[QsSٞԨ����XF�#��)�y��G���Ma���ש�4����BG����%egg_��	�t����fE���*�C�� k��SS����or.�{�5�|���8���?q095e��Dk���x]�m����*P]]]�[Z~;>KOO���?��	��y�/J�C-��[�1g�󡶝8U�`��e'I�4E��(I��}]�.kЪ����Oq�c���������g���܄�,'|��%���2�3<�}#��a��R_���I�e�n��8]0܊���ö����4�F����!��tK\�0p�c�$���;�6{�VqRRR ��3p+��!��aV����7���x%�ܾ//T�֠��l9����������DI�ﾗ��P�h�D��U~0��	�CiN���>�Ϟ��7R�#�G�q�#(�
-@��6���%�_o�Xw��w#@#�ۭ#�� �&�ߜ��ӧ�8O9e(N\ӫ_l�l�{�I�JL�	
����>B)�{�ȟ%UB�Sttt�L�&x�%�G�w���X����^���Ĥ%���Hg?��V]B�^(�SB�"�u[�P�4(	_&��q��m���y�'�4�|�٨u=K(T���qk1�W�WTW����l�t����*�Y>Q �.�C�UH$##���${�ZXI���n���v xП�g���L�d�����D�r�MοVF����KW����fT:?m�0c%�wCy] �RYYY&*l�R���;�f���#1���̟�]�ޗƱ�h��-�|�{j��x'z�����2|�ݏ��Xh���-d��_�Bxe�(�p��L
8���������;��ܗ��C���fD����k�
4?C�K��Im��`������ ������>-Ï��f��#X��#��#Lp��_[�� �9ӢJ4��� %lQ-�MY����lmm�Y7�%�m[ �CH�P�'����p�\O��7�8��A����=J��vz=v�ڀ��Qn�\M)��';r�$�BY,��Y̴��c/�eM{u=��r*S���/w%�x��?����'�x7hK�n�>�2c:���������a�γ��%�ł{�V���(����GAW;�}��̛��)��?#��g$Q�Q�|n�n1`�~�z�P|ͽ�vR��,�%y���4dd�:�y�}f�D��x�_����ujE������ �ml��s(F3܃�]�H�'�U��Eb������@���ݷ�2<�������2�t���i`��7b��jj6�d �]hb��8?o��uT9�2�7k1���"�$ l��E���4��A�\ �^&���g��_3"���?NA��q�6q.��]R$l�Ψԁf���1�0{v��^��<�صC:���$��E����u$7,�DB*�ŕ�S-
V�)���q���\�*JJJs+����Ϧ5:��%a1�YO��m,S�*c	��8�G
�&'S��_T�����!$�H�L��q���%��	�N�GB����p)���O��̀S�^U�HH����v-j�VvW�w��V�-��N��q�����*���<��O�4�i����ލ���e6">Y���3>����,�_}�6��i=;�7��o���e��t͢'M�qy8�2�Kmq�ts�Q|+���,��o��]��9���������`E	��)S�������A���f8X��&i��w�Xo+Y88 a������2)t�	���iz�z"
h���J�8݋&NB���� �>��Ihkk�XY���s�zG�o�o؞e��n�G���p�$䴸�N0�w�9�<��A��������l�T'��)L	�I�*k�����T�h1�l~���|�E7��ۭ��vE�kb��x���Nݦ-`���(�\Z����ص�Z�"*<͇�J%Q��لݗe߇B��a���Y�>44)B$6��0|\G.�0�R;ne�}i杚.(]���"z��Nf��5]r!�Bۢ�.�:��z u(����5�K��w^y��mU��N6�no{6Q�.�455���	_>��[���N��
U��4ݡ��ݠ���[r?�W�w�HGO�P6��~����X�n2Y��.뗗���T���a�.A�w0�CT��o��ıoQ�����e=�0x�����L��G�P�
Oۖ1�m��� 
:�A��EB� )D��0��ChBƱ���}?鿿o�#����6V��{�i�@0���_cY&� YH�"�������B=r(���;)����/�L�gb�zY7�� ���@�=�(N��D��d	Yل-�能=O��f��DW��_
0�Nǭɀ�m��s�W�,��,/M��ܙ_�B�����JV���1%�d�K����NNN�Bs�)�j�MTFR��ߣy����UWΣ"H�+���=�Mj�W�Qiؕ���|}���)-��ʂWՠ.���^�F��i�]�H�;	�3nkg�� 5b��EH�A�\��V�K?��H۵�H��v�~��q��?R��O��ښO�A��׹�����CUi�8�
�Λ��4����t�tCɛ������r)i���L��H�{�� o�|\q��?���~R��鋤��1������ mP/�H�T"��- G?5.g����q/෬��o � �7�!���%`�?�|�ص ;09�h����0�r�4-ㇶ\�M��IRz���Wl��I�?o�p�k�Cϗ�ME5��K�6��%��}�'??ߦ���ْ��"\�2 ��ޝ��&���t>]�ߦ)b������	���8w�]!*�@��Z�E)Z�equjG��0c>Z��%�C#��O£����B;Һ�3�{P�V�Jr[JU5́o�_�=�����Z��Tl�Eڃ'���*q�"+��pqe�{�F6z��{�Ώ6lk�����=�Q�����k����Vb�MǕ�A��̣e��E��M��2��W�,h�A�Wz���"o��������r����r19�R���
#�#��F�$���)4��vb��wE��1-G��*"*%g;�$Š����¯�Y����MW[:�ܨ�>�Z��9;m׮,f%Z�tq ��0y�:�ˋ}�����y��O��ƉaRT{֋��I��To�o�V/٧9�nF|����;����B�8�����x882	�����v([|Ѡ� c=QĽ��'�CK:���i�9?%�y廯�$�D�7%l��W��l�JH���|��J��8�	��@��x�C�;�<�>l��H�,-�^�k&j�����s0ʷ>���/���9���eb��U�(4�쥈o��a}+m}b����K�0�t��쭈ݐ�"�3�+,�sq���@v)����ާԠ;c�:��d��4H3}�D�Py�K~���ǒ �%j@�FR9�oN���7�F���COA�&�˗���n�~Q���ݘggg�mi��0+�zL4�,I������T�6��ۻ�U�[4�"k�/lY<�^��Yu_����hQX�SS �xr���%���%�D�F�mPJ�-Y}y�e�o�p����)�P<c�	Vub�ٴm{NQ�uA�)�;�-!8�@�8:��p�$��%6�R��A�~�����4a�"�p%�=�KO1�[�_^�ʃ�j�����9̞ˑ�䃽Nj㡬 �B��o����Es��v���,�$�������<|ͨ���r�Ho7>���3�Ϧ_z�st���ix�����Bs~q�	�S����5q+���3I�?��.��N�8�F#��Y>�v�.���ܗ�Ӣ�/��R�����1�E��Z �'�
�{T%���_���g� �U��w^��` � A�-Qd���1��/^VV6�L�TE�>��!��Nyp����c~~����;�>}z�*/-�sbf�S��$#�f/c����h�#��y׀�5�d	dt���7�����"���!X����.W�m�M�,�:�S�tg�z{:eȒa�{�=�^�v���2��Jwm��0�����X}�BA4��b"�F!�-�İx�
͇Vڳ��h$7X�Z�H��$����	
_�n)А��iEii�������fO>�����A�2B���kH�22 ж���8!��2�^(/�����5؈��<���r��z�\!&�]����<�*N�@5L5���[ �}�,�o�p�ma�p�糿�mDy/2���!�4����h'��k�����M��Ԧ�����!cQ�L���O|�$F;�1��"��Ux�Ɩv�B�c�@!�ЁZ����q���CY����s�Y�Cj9���Él:(�O��ѾM��e��&�������#���#��b���_���E�^��i_A)���.R�o��eNi�Pt�G<�aۖ��&+�XX���������^3) �L4_�)�)���#yj����!PDh؜�y!����>����Iv�R�Y���������g7w}Ij���[�=j�K�$%%e�E0�,�f=��:���񢍇"���w�Q��X}iXj�oj��NXL7� ;��X�p��f��k��7=���]�v(>��Y�Z���%������G��߭���Sp"	���ug5,�W��?m5�h�;C]d���<���ք4����|j~�^�5
<�qV
@�p�\#jIn�#/�o�H�cf0ڛC2��� Z�ߓ�	����U0���_�G�y��O��|��;�'nН�� ���6#bB�2�>�3���X>fw�]1tGV�)阮�h�f��Lh7W�vN���J������7�bUU����PQ������3����]�¯�=����ɩ�iN�����ᖌ_=w��ώz�"x�s�|H�VK���,>lły[�:>>��y4�����@�Aw��2��*�4��Iw��<̂��]=�,�9��{	�Y�w��{F.ݟ�4����`2qz�8���03������ʶ$X�b	z��:9R�_z@0�:!���������J��ŉ�j(	뺩�R̝s�C	|e)�h�~��pR(��İO�|���Y[[�΅��{�	��4�`t�����*�(�AU#*�K�n��������@����%��uP�|6�.��pVm)�ՠ��t�(x���h�\O3IĐ�e(9��C�L�ٳ����zL4��7��2I�l]E�嘛������y�|�.��\��A`�;�'g?n�����&�_����I�S$�̘������H�?j>��ʧ��HJJ2\=�g�a
Y搈��ʍ�MmS^7�J�����\���1o�"a�#y}�_�	2�_6�/#����E�[�?�.� V�����[I��`	eaa�p����ϛ����m�[�y�!��x|Z� 5���9[�X��:�,�?���3٠)��u�N�Z��\�T����2b A�����#���O���",�ۯ}�"�囤ǈY�jϏa�-�����͑<BQ�+m��O�	����9�#��2��Z���Ge��RC��Ň��O�	a��P�hG����vM''>��5GU�@��4�=qorZ�}������F�Gng��9N(��x������^���ǭIJ`��g�T1���[x ��t�R]8�"^<���n����w��Z����32���
���,|}�U�99BoǠ�.Cu_�kA#�IU�����qG,u����Wz�j�>&���*n�>?��s?�'3NK�^�K�R�tlӻ@��GH.=Е�I�&e�*-K��vz�=$�W�LO�M��WWb�y���b�-�)̈�B�=//Z?������I�m�$��` xi�P�oKvdm��t���	��qFH8�Uhݑ^и�Q��>����-��L%2�ĳp��´��N��]׆��⠹���b9�N���/��W;^�"n��I�Q�"BD��5�@'u^�* E�c^��ί&�É����h�z4l��m"��B����x��\JA�5�78XV�Vs���!�(�� $]j�NN:}Z%N������#�@�)'�����K+��|ݙ�����$x����������H�͜�}��oi����i�>�>R�����1���z?�(�>}Z��"�]]��뭭[D��L����@N���`��;�(������y�Ɔ�\+��.��2/v�T��BѤ�zT�O���fW�ݬ9fㄵ��v���0�D��3����qd�<P�o�݂U���L(�ʔ��*c�Ujg�z���v>$3�}30>��<4��O|Τ��9G�{DUU�`k�� �U|����p]]]åc��qi�n?ړ�8�[��qk�g$7��(��o��j1���>E\�ɿ	w����F2j�4�����m��3�
|�ۀ��"$��UҜ�|�HN�G;1��]�Md�����r냗��quS�������A�����?�z�/�W��5f@�ˁt'�x���t��"�0^�Ǳ&LGGG��ot�9������gr0�5�5;${�!�t9�˰)�&9�0�\%a42?»�w[;.no�D���ɹ�@GX�����ι�vk@��B��F5'08�ő�V����u�۲� ���B���PVx�[JY�?�s��'Wb�1�S�y'�e:96��ը��Ą��fƬ<��Y+��(&1t���]���CE���v���C�U(����ȝ跸o\��7�\����-/]�m��F����,�e���r�hp�Q�Д���;�e���}QN^?��5�@8�L�@gNȱ�}���l��eu+�2ʰ���{��.������n8 ��88-+��I���Όv�l�+9Е�ʖ��$��<� �d��0�$ۖ��c�S������h�[�y�H�vY9�S@�����N����k)�u011�fB��7�}�n���-b�zq@�z�d�k�~�^X�߆��{���3���H������%Y��]��F��[�K���fq�������%�KP2���E\����e1�f|+�E��Z���j���P��-�ׅ�������hDD(�I�1��@��a�3Zl�K����hd��-}F��'>���"f��(2j#�L�&�50�������œ�_�GHGY.�C~��}_���h�8,�+���N����^�#��P�YZ#��,�д�R�3�v�X{�N�q�?��:����^RS
�;r%����o��wN������h�M����7��_;ȗq�^��j�V����mya�`a���!C����Vj&@�fJ��\\\�O�˦�Cc� ��-��{vo�+��~w*�K9 ��v�۟��(�W���%��.�O%�dY����50@��C��E&�qq&!�A��=��gԮ�y[�8��AFQ�]�����	U�����60m�k(|4�b�G�����A�A<��r�X�/�j^�1��IH'^�C�O�z?c�,c�^"��cMF��,�j��)lQ��z?@�b|s}�a�͎T�� �m�)g8Lb�,���n��:vr�(�}�{����ô�,��G�"\\\�	O��
������L[��'� yi�K�A��@�?���6g�%b�x
��vw�m��\�㋧��bL���ݾ����8���0�	�ݽ�t�賷�3K���-88�#PeKFCC���A�Y��k���r5`sW2r��!%%�Z�����3u�Z�D|��w01[�^���}���v�NU��s�g��x�#T�;=��x��Atuue��58:�I�]=�H.
�-�W�E5u1�Kn�S�d����I���}���9���k���[�P�ޤ��>��t���ߕ���⿚���gb/v]�a��b��yh1`P�Y�^ ��T��ⶈ�-����ϊ�K��oZ�=�aZ��L��^V�e�Dz�/..ʷm	 ��j��m+�J�.Z���]_��+ t���Zz�|��ML^�y�|os�3�����,w��승��e���o���z�#����E�b|Ǆ�������Q�XG�`�7f��Wh�ubY���	X�3�4��;�O���g��pH5و�-�r�b�`����Ս��vR����>H����N�A8}_�aT�L>�'��SS�]Q��a����)�!4�VY!����y���!���ܴaY���]��Nn]]�ZF�fЗ,������7�]>Q`�	�<D�+;}~�İ�P(���N%y�5 �n'�@����d��})�x�]7
kNf�J?�5�^׾�~�Gמ�����9�x�S��T��o�]�l���d|w�^�$��*|&fy��tϞvQ~��1�PQm�ߣ^E�t��tHK��tw��t34("�)0�t� -94�1H����^���b����y�{�s�y}2�Z�ms�^0w4AHL�QUE���՚Wwl���P^^~�H-�r	�:D�R�@��|%N��� *�C���mS�����A�� ,�w��c2m�g�����N7o������ò���,�X����- �km8�y]�k�������gO�hi�#`[\���"b�7h럳y퍾��黗����-���+]]�]��m��M���{�j�����C�}+[��SY�Ι��Ϝ���?Zc,�y{X���޾x�S�Ë
�h�9U�n]��A�>�DVYYh�,��:w��=%���߿�G�0�@rlb��Ϳ�����5 gNc���������B�s�{{���(Y�����C1���!�9�A ��ɉK����^�5�Jo��#SS͓�o�i����P�1sy/+/���!bz�k�؊�/ݽ�}���+�Fl��:Ek@*���� J�}�*��$�mU��K{'��cQ�֢���P���.���&�i_�� �_g�4S
�X����8�����p�{6�^D�N�1<,,������T9�o�z��r����(����<���$���RUK�ᡡw��$��`C�J3�)��cJ�	H	ş6������f���'�H+���ΐ^^��rnT9�����".>����uyhwy#��5�'�[������E����_[X|���{�Uo�����b<��%�ՙ��O����:�i?>^�M3eѭ�!b}�P¾����nn�Y��L{���"�GR��4.�M���⟒�ƽ�IL7�n�EQ6,��UD���Zj��t���-����6==�ck���{P�۾��9Q;nF�	�l�k�P�qXO�N����TM�>0�:��Qu��!�����E�L�-����V�2���/�k>,�3�$�H�Y�����~���5/��ޞzn�{^<*����K���č�T_��s���b��5vx&hY�>B�t�+.�|q�V��M�vf����;�/�У�*�f¶&+iXYoC�\�����W�`�>�>�j�ƠH����L�i[]Rj�`�h��/Dd�G���'{�!���jñk�^�ץ�ͪ����;MF�.���i�RDf[*��(1�9�y��5)YY�������w�c�0G���`�۪�JRű�4�di_�t�	�c�&�֍���ަϦ_�2���X-c�ڵ��B�[�����}H��?0?"d#{���<��t���5�l��e:Il+�X��bt?��ܨ���^��Ds�L������)^W�c�_'���w���ձ�����m���J�û�%[:����+��'��̳���c�j�O}}E+lQ
t+��8��{��ʐJ��q�څ"�3��Уe/0gs{=���Vo�AbzM���'�A�7�����a^އ��R5ؠ�c��+���}��Y܅@�Ԕ^YEŋ�gK��!	�A ����nQ�n�xi|��8FT��F�_7	��L8��c��J��/x�}�d6�]&q�ٿU�|�u��U�@��b�M��BBcbbn���`����ҧgV8�(|�{��_�������>�.��Շ�����GBz{��j*O��F/�]�	�����������wo���ߡ�ލ��`O�DebbY
����*ъ������{s@��u�w�+�����;�僟��?Re���	^�q�q�|����e]���|��[���~,��IE��0���E�]S,���=22%MM���S�8�L[s[Ҋ�_(����.�����J���I����l��O�b�AmI()%TU�ǣX�@{ʐB�~�����z,229�7�u(��~�0(�le~&2侥p��!���5�k*/�$+�o*"?"���]!�	���WRQy�������@����?�L������z P��*r�Yŝ���T`0��m���bq�����̎�:���~q1�@+3�5������'�i���@�*')D�Bw����
J���n�m�����-�Px�py|�X�\d�;]!�$x���'C?�����b�p��5f2�D�b"�#�tX��]����e|�b�����pZ�f�(���T������0���3L�g�]�����a����ar�����Y�x�3Ӣ��ܰ�_O���qG��mZZ���p2�cE��U�U���Ó�r���	C_x�P�=RH��&6�R~��i�Y�:��ۯ�A$��~�9P,)H����L��k���]I��^��'5�	=�������X D6�x��s�Ҟ%��D:�ë)B��$$$�/T��-F��#�L�4R�!����Ѽ�������|5�)��}����1S�K��h>�/��H�����:d|��f�b>83�x�����̬��F:4��� ��P��Ʀ�� ���۫пTWk�џ��"��!2��t{�Q��J�b����?�9=�j��p�-��6KO�b��):�[��>z����N�	�Q���)?^1ʔ���XGd�KRWQy(�)���g�a`�ê�EnW��(r��*}F2)�`f1U0�4 �Px�i��[6�3m/��K��� t?�>Ya��E|��qq`�MMLXY�)���
��o���J�_�;iJR��ϋ��@h뛛jpxeMm���t!��iQ]]]uC�"��Ng��?8�rf�7�����unO�zɮ�WM�2��=��^"�N!�bd�|����k5��d�<�
I�6�IG��R�?��{�}]_��;Z���c5.V�
X�(D�����?��σ��l):�2�&T=ڪ� B��:!͈��щ�i�f���ɂ�\&W��^����{�]K��t0#��/2N��}�V�L||��r_��əut��
>S��n�1R@Df��%�0hV�1�?π���P�vS`����I�����3�Dyee��W�u3�܏|��f��[��Z�܀ݻۡЩ�D��z��icfb�Ty��q��9?~)�ٽq`���P��uī�_�|7�lϫ���q륳Z�9)���ۈP��3���o%m���h�iqj3R��Άݵ ���� |�����$+@��g8�Q���U�\����c��Qwy���Ht�{}�6H����=�Тmt��n{ز�P(�.�����	����\Κ/x�W����}��|���S�U/w�,��n5�Â�<2g�RI�w� ��ڢ��Q�����,����S���8��Xuʠ^�u�R16� �P�3o=Q��=rM;y�����%�s�s^h���h۞bim��\i��.;XP9�+B����%$$�^�����R�F�����bx������Q�� ��>����Us7��g�=���Ū�k
�D�����1.�'�Jj�SO�����y%�tU2j�;t9�t1FT��y��,���50��
Li�_����*�N�\dOT�V�U����Qt,7�7_d�󩇷����̶:;ܒ^�_��355�̼��������Q�����z�B"�����`xw�j�����8����쬈>E���.A�5����-:::��_��M�lUL���L��dq���	� �4u����N���>��� ��,��2 �QN}§E���!�Wa0�w$ab���V��=��L3����պ(��!}O�t2��|�B�z/�K�C�L����e�a�R��>-��3vm��Ѿ2{e���nO.��SR�r��!O�A�����bG�KQ>��2�x^�x<j���p&�,�n|�%v��5��~������1�7`�[0V0�d��?���������p�ә�m_g��$���A��q}�O�!��JJ�G=�{���F��0�tv�|u����E�g�k=|3e�t0�{��ޏ��N��x��/j��'�t0��'����EF��2>�%�3"���,�����$,�FX�7���JlW�����C��kF&iPV���ѽ��ֺ��Tac�}}o倴('G�ǧ!��i���#  ���V�o)�>�.�8N	 ��v)^")��8��ibAC@��	�E�;�a��O����q.��v�Aäʒe�sJ�d	���%���\�?�����8xr�.�]������B�3��p��j��{��-(Pם����ܗ��8X�L�m���C����Fn�֎�f\]�Eտ�Ю�����D�7�:�(�v=v�d�F~uS�~�_�A���#��uk��1M��L�n�:����u��c���[���܁$=
��;/[�c�n���a9Zk�iu>?v���yd�B�f[��4r�����OH(Z�Z�0s����w-/m�K��T��fi��g��B���k-��j����� 3���h=�VB�w�d$�П��/'^�M�IMY�ܛ����A ���y��+w`�!������1��|v^�l-��X�|ζN��Rٽ�d?��[���8"ǧ���<cI�O.�8hZʾ�O�����������8�S�?q2KI��x����fPV]C#(�������8�㜳+����t�e�v��K3J
���̽�~��4���4�IP����*I,�<��~�t5з�BT6�����=���@���V����Z��ޓ�1�ꇋ|�y_��j\��#���a��È~`"+l���$--=�{�ʽޠ@��y1����g�pD����?Ж�vSqʙ�V"�����>[B3*Η[Z�ǳĞ�0_."�ˏZ��HCӲN�Ҽ�@<��B�B�eD06:��lZ&��Hx�ǽ��
.3���aԢ�	�5� U��!1fă=��AR��E�S'�d�`j�����F���{p�����~��f��s��M��mo�m }�f_�߳ �Zk*/J�b�ު����?گ��[�S�����dt�K��r<��5�`�&IRRr�jtC��˴�N�Ѿ��~����v���~�}U�E䨺�s�H�xS�a��T�ZU^�
_x)tӻ��|T%éԹ��'U����+5q�$0�}o�b8W���E����x�S6$B=CV���L^�-��خt�:��\\\������+�i�2�HB���zD5�� ���֮��8c����%A�B�b��T"׈�q��UQh�c3ei�ങ�.0��r344�^w&����u���[-C?j�I�,���h����l�4�?�SQ_m^�K2Q�:�=����{��e�qT���,�_�S��l�:_��V�����(+ۺ>L�r#��b��(7W���jp���9�Cv�(zőhM8���!x7�M��`c��(� �[cq"��	�����[9p�/�R4A�Z��>�`cc/��`��%áU���Rpd�<��@��t�ϟr!� �¾]��槑|��5R����|�Y��3"�e[i����"r�yTJJ�z�������N���B`0�us,����g!��Mj��u<����̬����ю���d��OK+��AY���qk��`z�A\�W�9{N�����ard�i-��Vt8��n�N� {�xgAZ_PXX�˼7�s5:""M��^�v�s��KT�!.��s��}Qh=m����Eej	��-�2h��*�����:�ؕ� ��։Rs��-�,Mw	`�5�����F�b��9ԫ,y��Q��^}L��ᑑ��%.NNn�Sg���!��k���3u@5����K��4�󊺎�/,�̚b��QZ���^��;��D���oř'��Z�JUSU� s��ꏃ{M����A�ĕLp��5�M \�£Pb!�]?#���:�I�B6dע�5�l+A�������N�=#,¼��A?�U66�1�k����ׯ^����4F�t�0s�U�k�Si�TgPtq�w95��R%�*7�K��`�r�|m��`�o�*�Ǻ��4�@�� ��L��2�ܧ�a���B�Z�v"�S?Dϒ�T����_q���ZT�y�È��yy��3w����'�z0:�wO
�ԥhͲ�A��4ӟp��;���*]�׳PY��ny3j �A�DR=����2���b�V�ά�<M�e{zz�Q�"�� �.�=��	e���������y���DII	��e������xl��:�.vN�ݡ֐�9�T�Z�����r�=��ֻ,�_�f[=F[?������\K!v@d���A�/6ӝ2���,�N��H�wF����q0��Œ7C�ڴ��_P��=+�#B� ��u��Om+'A>���<v;金H�����>��|NN���p������D��X�O�<���◵>�g�P�{��Keoܓ,������ �����2�����gĒ�D�r=�y���t��f�[�ow�u �c(Һ࠮�~�u���y�=���hy٬�x>�>ܸ���Xj^Q���7R��R�(�{�vD�I���nQZL�X[1D�9�6���CJQQS[�T_�#xY�j��U�*��ط�MI8���vf�e���A�w�T���55:R�&��<�S�!��l��p^U�^ I���;B��{֠��]�'
�|��-�rt��"c��(�����I%���YY�No0/�Zit�1D!��zL~_�����[SuY\��~��o�㿠�y~�r[]_]URUU�v{����jXd�-J ����3d���üx�vi���ޏ��x/�^���Cft��}(d�����~3;�������ؖkO��'O��dD����K��9.Ɍo����᮹o�텹����&rY�=�]�5�R1��/	5]�ښ(/�����ߤ�;�tut|� �����؜��}FϪJKU=7(�Si�x �@2���C/�rS�}�vUs>\����ƕ,E
y���5�6�wȜ)����&�Y@h�yX�`.�D5�jj�����K��u�z�$����N�}���s� �0�M?wbbbz4Y9T���p�ָ5Yy4~�������Z9����65��VM��M��ܗ��l��SDX��+6��Z_=�/��ս$#��4k�^� vP����Q0�@iD��n��k�QT��H��ά��fo</��9��Kr;jٕ��v�Sm��A�4\�=�$4
c܄66�78���^���;[�~�J����\+1��2:g�ZE�l�,�� b�~ v��q�W��\Ӑ��&�O���2�'���5�F��Exb��E�Dk^�D{/7�}R8��i�ˬ�+���G�r_J����|�
��_C���G�h��(���Uy���K�%=W���A���P�[��:	��rtttL���6";n�p��5=���-��x������Q�=EB΄�5�c�2�,\`h���V|�D
��`�[񌞤d��C�I�@���@B��:n'J�	�*~��7'#ø�x��p�]mCԟ���>ꋤ(§� ���<���} {be �K�,����ͥ��O��.K.. ɏ?�$����B�x��v��})�{UZf�=����F__��):ķoJPw�nȯՐ$u�_��}��^�.Lx����#jY���U� Q�w[KA!L�*< Hs�����\}��V�h�H���3 ��%G�DH�7٧7Q�4�)3 #NI�K�FU�^	  h�nk{P�� �K�U��SPg��TPh*��g������٦5F��q4��+)��X��+>�H�prR��yfhiiY��t;0J/^����6b�j3��H���[c�'�T�Sa�ڌ�n����F2,SY;�՛�������c��G�EbAx�������E��G�	�����n�k�R�ɶ���]���;����%�W�-�ٽk� �rۿ�CFc_l)�N�c�����VJ ��|���<�8��x��X rCc��0˂IXUr���x��]�;rM}m%%�<�����i���� ��F p������Gp�4�q�����qk^��FQ4�`�9��c�t����eW�)��\���4�=��������^;��-J2��:{{G$��3�8-k�,N#��>G���.��Q�;BiM�����+Ip&��}4�5I 0,
�a�ĵ�mw�j�N�ҵVb�! �S잩���7�[��-����-d1Y��Æ�wRt�
}��D����C�QZ����~7��%��z��u�GR�j=07�zB��i�	���	��6�@{�S0�+������S
�gׁ���t�+��� ��z�����݄�ֆzѠ��j!t ��J�a/���VZ�L��o`�7�8���y�v���[A&>q�6�����v���٣3�CkDg���N&"2���aecA�d8��^�S�ˌٷ�����-�@|��0T{������`W2
t+m������j� Z����${o#��}��ؗ�YH��#G���������K����(�S̷�v�Y_2k㌝EL�#��K�z�O��#_���q��s3"���=��Q%$$��K�[+#rbl�v!���?Œ�Z��� cRR�z�R_��XbN�\�쬬TMM���h��R~C�*�'�����#�T���wD/r�C;���-�$C���LC#����T'WAWn��/u7hե�%::���켭�.�#M������Z�����Ɨ�>==>�8<t������5��,���-u�hE���M�iM���_��c^� 1��UK��v���9iii3^ �+�fD�b��u���F߯�X:�O�)����		y ����"��[!��}ް�4m{�ڤ�+��եK똾���o�n}o��p�f�rFH@���AZ 8 ��0�����WN9���6l�w�^G�e����o\��5�I�9>�S��8L�j�(��%#'g��Ǒҗ��K�s[D�7�h4O:���|+��|�Mӓ�n�R0M �V����7:�S��}�i$F�ݻ�����hsH�RO�7j�)HN���NJѴrf���
�tI��VE'�K���:�[{%�*�6	�@�#��\����tx�v����ABX�+ /� �Xn�������W��MWw7y��́���K����S�:U�i>|�2��q�vY��d �	J�١�8Q{�cg��<�^�w�`
vP"\,�\[8>���90��rn�j5��?�B�A�5'�	��VOy6쳽A�t)��K��Hŵ���ƍk�ӌ��,���?�� �G���$u���|���		�	=f.��9�U���dCkKk�lfaaaF+pi�f��O�nYO�XK)3�K~�����X��`�]�
�ݿ������N���)��vϫ��L �y�K�T�f �f1RVMI�������۫����Ѫ�/�$Z���ā�j�ۓ���(6���QI�~�۲��)l5�BHDԵ�Ki�8���q:5�2!��
�9Fn}�������Oe���{�򤴷����oa�0�M���4HĻ�D�,��J�EdgK��Q"o�M�@�6ۺ���q���=$��~�PLK����n<.F�"7��~=�5V,rF5@,0�e��茢g&�F i�%�h}h�`¯���$�L$����i���O�����g��q�pV��FY�������F�G��'l>�s��	d�ff���7a���� ������6b\�/��:) ����A�.窥ބtt��-~̒�Jl.ϖ��jq���p�)aI��ǔBnJ�L���(�]Qu���76]Ӑ�����n����0�1��5�8Ӧ�Y`��D������ţ3S����'x=_�A��BTԿ���:bV%ElF]�s#�j�5z��Hi���ϯ+��0^tI��Q		V6��2j���>�r`����m5��t*�A|?���<W�㓬Ivs�b��p�����]��)vrV2�<��u>����9����,yU��3��j�oo7M�P��
 ���5����tx�� 
�ܽ���Y���8�yu����W IݡFsQ�Yڷ^��,���3�����(d^ƕ���L�s d}s�3-��9{�Dl�'&H��!A� KOn[�:�<���2z�`D�y!G�.�ͧ�M���P�'<Y�W���Yz��ḣ"O�2�Q6@���*�,���j�m5
}e�a��􁜇R�3��Zvw��d[[5v���8n��&(*�i�ϗ��>����-(����=�Ȯ=��?+ʝ)�z��/�U�.���O0>�����������@���: 2�9dѣ�s���������>�h��s�Ky�+/&>�����}~|V��{.�Є���S��u-:�S��]7!IRe�p �>R�X�3'}�%<�m\�9���H*#UV�o+�����Ԣ
+*x����p��}/={� ;��A�\ �>��F�2�H�����/�?��׊"�I"i��R_Hb�7�'�ܻ�ڝ�p�#4J����N�cWggg�	{����e���������"Fۿ�aMW]k��F򕽽���AM^���a�{�R:�Ž�	b�Dh�IIyϊ4؅Od����X�qa��
�˃1�!Jx�����D�iP�*�"�C_��*oMU���ʦ��7�����S�!��r��$�@�A��U-����Tp}0�OcS+j��ؾ��K�����-��b�o��I�"{�}�f�;��4�H�:�ѭ���*q�G�H�9�(�8;g�?�������u+��A�o�aݟ��[�W|XF���_K�t>S�$�Q]kC��j�<�l0��~ ��;�Jߣ�T�o-�;C����� ���M&|^�����3E�!_L_����Ȭ��޵��3����� �	�F%���{�Û�t�q!���3c���*������TZ:��br>0��*$���'�5Y���~���B�$�YY��P`3i�^vE�Idu[�D��#5r��k٩bX��x艉�Wآr��c���xЫ��	 q�+��WZ�Կ m�Qy>�j���y$�&�c����i�����cia���ނ�����GAZh�=���_c��ۍ�Е��7�/Z�:�D�yc���I���E5�bW���Q����	=s5"Y�D������JVV��.�� .�0F��,��Lq� ����Q�B�F�"0�����S����7Pl�b-9`$u����^7O�uM​|��6.d�!�֮ϡ�&{!3�[*}y����N���5w.`��2i����d� ��3�Ʉ���lR�[o��H�h���0ųw�{�	B��_P "Ƅ�,%�`�,�<J���S��4P4��xI(��7��M8���:зu�2E���_�Շ%��B9�#E�#H~�k�d}��m3^"�N��"�7���v����cK���)��hI�0���u'���y�eHT�<�k�����s�@�3H;֢���JD��6X�9P�1��������Yr���T�!�ا��HP��0pX���^fg���D�o�&x���}�!�0���n:��Nni)W�4������S�w�9���2TVN۾\�>=ASU۝��$x���&(0M�4��my�8~��,��	O�(=}��8�/�5��`�����T���dh{8�#P)�.�Ϟ�>�b�60[��9%}�7^ة���f�wk�^t���o�ɭ����_xm&2�@ ���YH���T�u_*k3�c6{�"� N��9�ū�/��)L�yX]Q^��/H����)J�Q�m��d�l$4���B�o�0�����v@��X���Tl\⟝<b�|�:X� XvᛂTǡG��9�/���>J��N2QY;c��ۇF��r��մ�)H�����t���0t���Z�hYG�2�&$+���M��
�Š̑���,�zyX0�W@蔘@��
��К�j��A� � W@z�["�Z�T��ߣ=�q����{�	ч�{���{���4�7Q%*�b�IxA4�"�FF4�s�iiϊ�����rsk�}��zUL�s�IWYjV}�����$��vǰF��)��g�(�-��_��i�	-AC
�p�z�=���S�s�0ڜ�
CT�Eʞ��ѳ�8>�m�g>,!
w�X�+�ĺ,�R(H�T���K��L\\Q���U��+߾}�%1�i0f���j)�O�b/��.^vX "z��z�G��ƛ�l����ut&,����FN���@�Y_ޏK��,��KnII�Gc,�J�'U]����x����<A�x��e�篫�\��-M`���e*��D"��F@g�tttLH������`G~�y�F��L�'���^s,�������"cZ�e�ju���U%]��{��`���������:���x�h=Jg���i<I$�r�mmmh�٪�O�4گ��� ��8)ѪhI��7��Ocמ��ר5�O��uY{I�d���Sީ:Fҋ}!�EEM@o�5�9�  Y�i���J>K���S Yy�i]}��03E���^!r09�}��*\-�y-��q##�.E�F�MI���J���~�F���L6��^�aܔS�-/c?�}+�����y~���2a�qE�;�#�FU�Ⱥ��^!���?�M��F��`x]*#��K�A+9R��B�U�ooeA��\<S@%i�����.>+��h��k��Dԧ՟S�QK?{T3��2�X;g�HN��\<��^W�JSV'T�_���p��,���摁�B�!�ȏ����5�.>���qlM����#��n�_*�xSQ��p���d��W��-7Y4���~�� <Qa� m9R�xi�ie5QB=����=�t��qEQ�
�<�B o7nn�i+=�p�ǣ��{��%`U��,��ɩ�������z����99��q�̼{�i`�&�x,��%Pa9 ������)p���u��n-��w�f��Wp��o/�}� �V�,��Q!�������-RWI����q߰��p�F�%�|i�-�9����8<��o�|[q��Ϣ���*Tߓc
�}�ػjN�P)���E1̔��F���]9�E&�����O�������sO;�8��V,.�Ɵt1l��3:�K3�R����ɖۡ�7W|DAa�OV�1u��x�E_�(���f����Z�^��,��8/~
�؊�X���9�Ġ����& $�F��vAF5<ϴ������_��'_5�WiF��>l�f�R�
t���I�V��F	/ԇ!PK���E�)���^�0�����a�xL׊�[�����t۪A��[�#!~�
k*��v�������g�
����������q<Y���-t�4y�cqU����QjT���F�<���d-Z�=�Vn<�x^.��<�۷�G7���(N�q������W`^������������*�Y����Mӎnvb��K�n��\��p]&'���}�<6�w��~��b6����[��С\�)�zQr=^��i���u�)����ٓ{/[���sF�	�4��q�D�a�g�����B��h�Bo�[�����tOQM�7x�k\��?ȷ�T�r�/S�Mci���D/��O��,���TF�O��%�E=ă�h�6L���d1Ԝ����_rl�?%�G�P1�����0���|Ի.!�/���T߽���NE��rnx�L�ѓwm�*�o���G>ky��)��GK��Ѿ+��|��|h����p�BLJ���e ���b�xH~ԗT4ި�����C�a�����щ7�MD\�����Ş�3���'m��%@�dw��
�~4?;rܮ�F�R�kʊ���4��O<]�Ϲ4e�47��k+��3�{◷T�I�%�]��N Z`�Ģ��;�\�ܝ�����_'勐b�f ��Ζ���B�P�������5*2nM����Z��Ջ'�-[d�5�q�w,�w9��]5�������-�O��IU�kuH3�C�����\$9�v��t�>��oJYHL�l�"b7�N6m��G"��>�[۱ިK�w���I�,2ol�E�#���.�L�,��Z�P��&�r~�^4����T꩹O�~9E�v����hQF4	㌛�d�^����������*��Խ<[sԈ�M��n�4)c�..��{�L���h��0q�����P\+���QDQ�&��x�5�.���Y-h�� ;�m}��f5hǄŰA���R�_FV6�F����-�@������|h+h�8\���=J�q���"[b��wu�>+(�y�`jS~7������2Ʈ�b}���@iT;��ڎI���@������8�@��!?��E�lc-�����v�+�� �G��u����3����*�rrh5��Q��b�G�{FK�F ��5�=�^.4�5��v���x��p�?��يHyݷ5
���!���-i��J�Y�ᮺ�	.�X����;m�<kv��:]���`X>�i~���Fo�%���9�7����{Im�f1����پџq{�6��|��tG��X���>���e�p�w�Wm��4+�QA��F<�I��黼�u�lY#|��2�\�s4�B����CR����8�󵊟D���'���@oprr��l�������Q�F�i��uB�\��w+�S�^7+�4+T�~�UT�n-����m���zd���	�MK��*����kI���_�9;ʫK��	N�?qZJ8s�S(,���'XK\�Er�7��4p���~�ν�0����Q=��C���p����O�B���������	��l�������$Һ?�κ߳�=�dX:X?��fo��Ϫp�M'����΅Rqm?���Tg�s̟��䚴�ғ'�����3��FE�fq#O�U9�ߓfii���2�m����ѿ��t�	���#����H��߹nOD3kZ��&�4x=�������7�m��:ar�O��	��Jzq�V��.�����+�V�T���*TO.Umu'��x�k�NDZ舠auP)VfV޴�����b�tW��Ek� �m�g.��ae���B�<���;���ThƸ�:�m��K��2��~[g.k^R� ����n�̅���i�{�[�b����5kSD&qU�X]���-�X~����QY�yk���v��X�ڔXM?jŤ+�(&��L|l���.�_:yF%���f/u��ed�����i[�7`�s�$�91��}�B����Y���bA��d�4��(Ң4?��UHd��q��!=�u[��9����.AZ�i�.�
:Z��H*"kwqA �$s������<�@��%�hϹ�Ȟǖ8X�р��������tSh}�X'�1���\LVz��q/f�*������f.��v��.6�o���(ۺ|�� *6�>wZ֦�D<<�������<����"������M����b_B�(�ͽy�#A@+�����6F@$߾)����1���!L$�(q$(d�"�PV�6��h�(o�(m5Dn��p+���񝳥��n;gf��ُ�V|�GgKGg�11YO��o�ao�Zd�!%�����0���U��������ޜ��wbI�yH\�������n��dVi��>�X螃�GMJC�G]��q���s.&����b~p���@s��@M]��z�GaV}d�Y�\x���$o#��r����".kw[+o��"wX:�pW�j�L�$� �sO}�y~��օ v�=<H�`�Z�����	�\���w�j=�;�0؍R�Q6��FA8zh�5�`HU�e�m��ܪ�L��aQ:Y���ҎKr�2��ۑ�T�d�8�L#��nA���Z=����݊h�������Pf|���N(M�i�F�Wi]�g}q��Ӥ�'rΫ���Ӣ����[���C�Q����(��Nu(�|�D�$��w���S��6"���{#�fa��G�9��E� �tv�:{�H&���'��G���Q3�։���H5���Ԩ;�!m3���k��}�j{cᄅY���?<=�WٷU���5$� �m�KJ`z�=`*̸)Y����Ma����?F���G��XT
"9p�C���$�]� ٰ�ϟpb�S��%
'��7��	�_}%��'l�^^Ssk������A�xu����^;��S��'p��z��z#�W�qB���
<)uR�tø�JQ4�cwa�ɖ8m::�]�r�H��f�F�H����;��D��^��)�t&��ݲk�z.8�%�]����ؼ��~���rK��B$m�	Nf��=�)�ō��ڢ�U�~���9��G�?�h�Qn7��+٘�!֩��!fS�@�<�>���>t�&`~o�34=m���4�V� V7���Ą%�E�ʫw���fc��f�T�0*e��P��5��[��8-��"}�]�B�rt����l6 ��5�gd	�G�q_p
����=��y����(�ء�J�5>�]n��g1pc����z�<Z��i߶�Yf�F��9�.��g�Mn+�HuP������Q��~��_3�;���@F7嘑B�3��Y+'YGfv��~]��n�W�{\.lsy�y���+޴��%��)M�F;Ĝj�r3�(w�<�1�^)��w��M���k�W��}F%my�fc.�7It%�����<��3{�zz�k��Kx�ޓ�C�A��V#,�)�	�Q��Y�;��A@���J�k����EM�ՎX�r�ϒwcԘ�-�Z�@�O�zN}}���
�Fy8�ܝp<)�qqz�W)�Rʄ'��941�����=L3�j�����(�0^rv����8��,����<�Nh��:�@�><2�%|4�t������z��m%Q�75q���k������%�K�(>�i�t��6�����Z�-�I6le($�RԸlT:5`��$�y14LW3����zŊ����Jzs�!�ڭ��i�k`�4 @C�ׄ�F�q-ɼ���T������L���B'���SY�%�m��yT	_'��6v@�~2��=�f��b�j�{�_K�v�D��<�:��y�$?�A��X�6P���;S�V*�mO��u%�9;�
��K$eM �'���\�Q�Rq���8����q�[��N�R��C�^���	�er�6����씌����^љ�
SM�!�p��$�����i��g����7���su5�Lh��`�ϋNsl�`ª��*|c�rfDApˤ:O����G����':;�ٙ��qw�"+B�Er�����l`1>�D&�G?��K��ύ"f��^T��7^̳�Ч�+cm�1�����@�>��?q�u�վvsӊT30����O��c�ׯ---����i �w|��P�bb��7BP˲�佩�.�&����0@F����<,*�\*��x(s`(,�+a��{A�i��0�?#c£��feC��t�%9��� ^�U�p�����N�F����K��]�G	�Ppߘz�Pu.�=ԧ��!L�AX=��6^�b<�o��6UC0Hݣ�]7��X�M]��t��QM���^�n����[�(��n�cY����.���?���׵�BB�%CGG����ոl�JC;�S�N�+�p�ɯ�����[_U�}=���ȃ�(-(�-�"�%����AH7��0�H�Ѓ"9
�C��Đ��{/�|>��{�Aa���9k���>�И#7>j��?��.�V��=���@g��U%,����
�s�o=�l��0ඞ~Y��>'U�褨��L�:&��A&��UC����AP�ZOk�����W���g< 9`�ed�(2�2�a�;|͹�3�2kR��P�S�:X�r��Dl%`�� v��`l�&�����%���J�����rUK�I؅��y8���$n�g��<�V7Z���sO�������b�`ss�>oRhh���Ժ�q\�:���J���n�Ql���K^1�؟�V=F�+�iVr#1���ʅ.|�g:Bŗݰ�\�I+6[S)���,Ze[�@�����L��2�q�2��N��RF�?h�]��!!%����N
C
��t����j���`��� �9|i�+%��:��<�~q���̜x���]uaf�4�}��~��^�R]�~{0�E]7U�[&�cW���
�=#{�� ���S�/Ow��'���M�#��E5r��%z�m�o�7|����{J^y�}j��2";<���g!�5Ri����B�]����5�~�}�w���`�S��j�$@��5d�N\�}���u2�!���r�c.�$�M�,*��=Kj��Y��N������8�C���S�C�$�_|���|[�;�u |�~\�y5"͛&E@.kD��� ���et�qԧ���8�<�*��4��.�9-��O_n�^����꼈�'sz�T�7���(�u@�n���G&C�����GT����4�gw�(|:(�h�E�D�Z��ݨ���'��,U�+b��˵�P7a�}^��Z�Vg3�f�,K�/��>:$��0]_A 봰���3�L���q��?&ߪvb�}�%iDdd��v��v20������%�G���ڧ�{��8�$�VM2�Տ*@�p����$�kFs�cE_pl��z��ʮ�Z/q��M����n�~Lkh�_���7#���6_�L3�3���_�9Û⺖�^g�y\<�1J�ȱ�͚R���ðE��5�3O�#��	�S8�;�ni,f:T���nj���F�տ���mY�n��0�}
�EdPp�H#P?U��X1+	��Nj�o����J��!l1��G�O�^�[w-q떦 �p���C���eB ��k2|����\'�`�b��Oma7?�IS1n?��z��Z;�L	�����W�:��Z!;������N܀���g�`�y'3@&�]�Ε�|�п� [l�X���I!޵ۢ8# �q#���yPD����PR�l��A�]�g ���CCZ��)���V��b�(�ɾQ;�z��Ip�N�J27	����P�� ��ܝ�\���[�C]�>��Đ��~Q�%OѲz#]O"��]#�O��4�Ҭ����8���Xvd��9|�raŜ<@7uT��� ��IQe �"@��^^�xߗ߷���Fl�[d��Ie��k;���}4\��/#��'XR)~ݎ#����� ��K�$���glq�����)s��O�&&&���K��	�G�R����u$}�>�����G�Ć�jg/��b�Y����tjO~4��L��2�S̘������A��c���_9칠W4w���V)N��G*��af��oyj�~���� >��lDo/y��)��dʵR\�=�RNt��S\7��4(Gyf0Q�s��g����n��ٚ�(�i:���v4�qN�0�4��|&6�@L�=ܿ��%r.p䤅@�6v�l\]5�̿�3 ��?�8�չ��;X���^dw�Q�)y�o���=HF�����#|�轸h�[4�fu,��;L��FdB�^��&<�e4(�n�E��T��EJ�3y�����# ���	��w�_3�9�so�DTFXd,�}���ƆNwe�x�%�t�O2�Q���ۮ+?
��M�aDf v;x5ZeE{���=w �xxx ��5g�lp���9�aT� ��M�RQI�Ƈ�r�}����7�u�R��&���C#��)�7A�9�k8� �a㠹޲��m��4I����Su+>a�+3�kʽlɤ����JTt�Nf�0f�-Y��u�bK�a-����UD��
�;��#�Zr�Up�wD��\�D�Y��	S&��,�(U%D����p@2!z���ľ�B�C��x�/]b�֙��j���(#�r;��W�Z��@���1)��<�`�/xGE�߈`O~N�K�Dc�t�h�x�E�J�s��R@���i��n}<�5ģ���"õD�����3�����P�- ��e>�]ls�	�.�+K�5����E~�;�OX����{�%3k4g��!p��Ps�)ǶZk=�����㗤�v$?�"�Q�V�؛rz:y�I���~|��2�W�1�@I����k�"韪P1U<"��>�}߀Td��!��PתN��W�K�F5�1׈*���Pϣ	���EΨ˴�g!�z;J�;�-k��r����dU�v:2U.�ƺ����q	�?D_N�����}A�{ඉɳ�������a��A�A���6����ڟ��7�:^?�lO�T�@�S3Pǚ�|?�^i����.H���z��d�����Tw��;Q�ŖVyt�ȸ�tP��Bz�d��Dl��)b`�iw;�{Q��G�f���UM��nXj]�b�З��dk�I��Y]���X�ks��O����pǖ���7�j�m99� /�ėS��---�� [f�bn;Z%||��Ѝ�x�çCO>U.t`=���<�F�|M��ښi�ҡ�.d���?�҆��r�=�2y�2�+��L:��������Z޺ő"��!�}M��a��\i߱��8n#q�><�����$mjMu��5��]�$�1���z�ćq�~���^Z̿4~7"�����jx/N|�O7ZK��[g�s��=WRx���q�ed�Qo��ۄ[�u���x	ֽ�0PY�ٷ.bT"u+G��`���D&���j�2l|�hT#��s$����l�&��n���T��\����&���K�<������{�������5�nV�17R��A�L�|<��B�y����(Z[\��R��QJB���TRf�6h#>M��mi
v�M2;褋�ܢ��``�A�� 4t�^׻��b�_�6j��q//�-A�M�M��^a�!֪e�3��hh�1���"9J�3��,��7G�R@Gbt,�p�?x�B"�v��Fs��b����G���'����{[�a5OM��1)D���C7KLHh���Sg�T����&�5u'���E���1�����5vI8ť`KK����% \��{#����x��C1�4�����x4z���zc[�J��~dmii�u��ש���*M�[��JѸ��Eqkj�P��Ƀ��x�&nX@2"��p��(._߷�Fjw�� �}�*�3�#�S����5�[��m��ʖ�t/#dc�9u¬7�&��oqKz�X��w�Bۂ��z��� �?�D�ή\ Q��[�9e�U;��η�u�4�T7�aM��9�rU��ر��5g%P�.R�'�|��^���ѡ2��w �^�C�e3*��j�˔�S���V�U����_.�U��sN�zԑ�z�V]�S��sLT4)|Qg<��B�^�l}��y}#ڛ��mGh1��2id���;u2Bϗ.o�Tm�Ib�JJ��ڕ|J�GT�{���z����������_J�#x>08D�����;�~�n�M�$���G�k�I]�S%r��fOn��z��=-��M�s}��娗�]��=Z��#�GmuU%���Q����&]��8��I�@T�;a�i<����K^z#?.�0�S]��/���}��y#���qv���ٝ
V���Vz��då��7@V� 4Fu��)vx/  �՚��������u�%p���V?��u����.���(&��Μ��"������<���ª=Аd�=��[i�j�#/��^��ʅ��;c�@�s���%���d@=��6���S�_��nY/K@/���l�N���s+�*Y*-�l=��H`0��;b_$Ѭ(??hb�Dg&�a��r�mx�PE�7��R�
�7r1>E���LS�q\����.[���5�ky�\��3�����S�X�.�i������V�}j�������'��}S�^��K� �#*d���,���+w��̼E :ⓒ�����k1�����i��'�!��J\�q���k�5�7��:>�\����Fb'v�Vq�p_��y��\c^����閯�K4t���"��V����]F^G>����Ѵ��\�jc�8����������@d�9��V\�~��K�Iۙ;:6���+�v�d��~f�n�P��>*��F�bg��m{��o���q�S�ҳg�9X�ӽ�/\*��g*fϥw<27�G�7���!-���j��M7�^g}*�wP/A�h!
��s-�c�slʕ���1�=`����L_�tp�p�
�_���1k�X����B��&�e��'H�[��y&G T�Ҧ_� �a�ت"A��g2�mX�&o�u�n�����
yq��V�!�x�Y]�'���վ0��a���Q�ҧm�]�	�[��2P��Z"S6t���<��(��@������k����)����͒fyYG�79�� :"���%(e���j��6W�V��A�"[d���?��oj�0�Km�]tlU$ѡ �N���(�bά�;2!l�Ud�l�(���֕ ua�| 5.�� ��s�X��`S*!����������}��H��0=�13��������C���^�0�C��v	�MrLj+��@���w݉���7b&sy�Nt���6I�x�v^DB�A��]��zn���L[�����с5��7��ߊfe8�Zl����g3��O(`�V�)�$(͙7&h�$��j�W��nha`��yO����t����S_�N|N������S��z\���������{���-F�y�b;�� �����P%�4 �[��A>��n1׊�x-�5�N�m��r����Je5ӹ�H�-��.r��Ƀ9�|-UzSe'�����Н�޾=��pP���<"�Xa ���f98|�2�(�`��}¥�ձb��ҍz
(��ru��$�Tu����L��"�Nxnܮ���H���	~o����q���I�u��D�F=�"���-�:�R)h����;zU�w,���l.>C�Wk����wu�@���`�'&V��$�'� �z�4����5;�E�"G7Cͼ	?�9(o8��k�T$�aTE�I���1��7ʫ�6�}4+Zn���9��1��`�;�i^)=�׈���E=~l�Z�@�^�߅4W�:d��G�}+ڬh-��N&� =�v��%s�.��Q��(�#�a�RՁ#>�b�f�s�z�FR���F�	��d��.�)hT�A:�(�bI���W��Ρ��{(**ඬ�/ "���PB���g�U6m�'�&�9pI���r�[�zJmq
�'G��B��̹�F��OrK�W����FB�\�sT�'\�q�-7��4�?��7����c��/�9�=�����h���^+�; �bCC��c{���B�VVW�W��^��V�i�P�5������Q!b��ˠ�ܠ��12x۵'���*ȏw�׭ݤ���Xm��\KO���x���p��B]ʊFG)8[�њ��WA�w｢'�!_�,ڥ�^�V|�v(���ϯ n����-��%�/tV�s�`:E�'��Nm��W^�b��ҥ�����h5����x��|.�j�{ls�V���!S���'Ԥ�ٳ���]����'W����\�.ߗ��4��kZ?C�<�}X���MT�F<k��Yt``��8P �MLL8��S�*j��4���SC�����˕kz#���p���E �0��FT���l�����+�Ic���?�*���a�E;=8J����gAH�҃���݊ļ�(�b��ɷ��n8����P��T��B���<<�b�~(%�%��3�^R��B���3|h������X*��o�׊ �pj%%}��n����0�'��{�k��=ș��D���Bod���Q��Z��L5W|��������P�j�6�CV��'7xF0�cG&�23f�<5�c\w'�@n�3-ND����s���8��F�X��!g��Q�ŵX5M��R|8�S&#k!_II�]����0#���#b�����Ĝ���q��cH�f_I�:2agP��#[��^�9�=2n>W��j�,L�D���稰���:��VC��+Z;�O�%(����ï���{� n}�N���·Cte}�F0Ӂɵ���E�=k@hٙ��������@�`�C����I~�%bZ	�De5�ӳp��j;1�#ur`��)E ���|fR�B�¢����"D7ٛv��G�����f
� ����e�շě�wҬʥ3�h���|�����^ʥ�8�A�Ѧ��K#��.�g��������Z��w�{�����:�l~3Dc���Ԫ�����?ٳRϗ|�0>�^�f�3�^%,�6{Eo%l���5�3������O�b�Xk;;�S=��s��s���zj�Z,��z�v�"r���G�����n�wq
�C<W�B���c��u��H%3i6bHmr-�3�m�j	X�?��4}kB�M��Հ����6�\c���G(�3�A�	����`ُ�0}B��ڌ�ho�^�z@�W�׵җhO��c��g0���>t�3����=�o��ɹ�fn�iTL��ߝ�N���Jn���@ �#p���<�h���Jm'�oǮ4:�X|S���C������iy�Ў�]]mP���!OMF�t��?s����+.=���uB%����:���, 1BY����q�c*=m�M����,G�j�[d���z>-�-��]�\]�3<���񛝀���rmWE_�Z?5Po���%ʷ9�j|6��|��"��ѽ]�z�^P�/����q�x�2kTB}��!��	�H�h�=�b<�Gc'�'2�z�~0�;�0����[���Mm+e�{�u�f�U.=��+;⻟�%2�	8��+++�{~v�2@�u��QO9eU�4e���-�==�6� bv���0�����V�٣2���1`���3i��#H�!���4�Z���6�(����)�֤߽�8���8A2~��~�j�o$<����81FJ:���^"���[kT�����,�����E$hr��A����% 5nL�*$���L�,!G�V��XD:��F썍��6��IW8�Ӣ�H�AB�]�- ��&�Rg��6�0��z�s�M�z����w*.�sk7WD*��t��Qd� }����ȗ��_��H��G�+���׈��@���0��޳�<������j.6]��M_gg��.�����|�ӵ~{��/�ܖ�"*ʌ�V��E!��m���-�7�O��w�&�4܆U�p�0Z��� <�ke�>�i	�,�[��gkF�qRd��]��چw����]�_
lq��90����J�=0^�����^@l�:B���_���a�ɞY�n�Z�"�Z��3��Cm��/����C��
[3��ː���MO��M{{U�O��|3}�t�n �8c�՛�eUo0eB�t��d�NK��A��]�֤�&�1g�x�>��Z@��"�`�hgUT�����Dúz���p`xi@["$(��6i�+)q-��3���;w� Ln���+/�Y��I���{��r��H��5��C<=�Yf&��Z�ͬ�%��{4Wp/��6ƽ�������$Da��a��IBc����5�h������^/O:%R����I`�j���֜��zz�5=9����[2��l��=̔�c���l����d�}�#.�x[`���>P�Ga�l_�#S ����9�
��G�{�*��`E���x�^լgO �	��������nb�Զ��Fм
�f���dԫ�	��Y��"��G�Ɋz���$�Dtj�w�uw�k%�� 3:d���Vy6]�f$�/���o�J$%� )S9��}1((��i�$��߯�t��=�2�XGG^ri;M߬O����[n��a�LTe||�`��zQ���(�S@)� �4��v��Z�u�����'�ydJ���4I��I���1�>{(T���H����q��x��Un_���Mne	�M�k@A��8E�/I�~x�C}>{�,�m��"�X���B<�29(�>@N~~<2y�o��^{e�(||`o_���K�ug?�oT����oHO�	� ��D���iNe�c�`��vuբN�����z��nKG��#M�Բ7"�|�.���t��]g��3؞5�
E��|!#	���ۼS����_s�@r/V&���ܰM����p�u���#+7�՞�(X�`[�㜉�	@�f��!v���q䌺������ވs�=�l�<��5}��Z���'^��6l@�ӏ�ٰk�HX��TT+�x&��Qw����RS���2w�b?�d*�.Հ�Cl��-Y2�{36(��Mzz�?5ï�u$O�[o#� ��� 7Y$z�:6��5P��i��5J
�>���%�
�9I�y�bk �}RNh�G��l4��:��R��e��C/���Pq_p�����i?�����Yu�
T)r9�zl���� נ��������biY�#�UX��R붇���A���D���3򦍒���@���I��X���-+Fߋ2m�/I�U�=��	� ����	���?�r"Nkg�0�Y���l�qR�<�{�%�&oU�f72���Δj�*��* �^8�+����}'e��R<ڮH�ۻ�c��Ѕ��l�ł���o�īh�Ǖ�h���Aq��_�4���r���X�;G�\�v�X+�n�}�$��84
vY��1&X{�t�@�R�!�����~QvK��-����h
�=���C���@K��FPJ�<���BZ׮��_��O��Yԓ�k��c����n֌:4=��hd�O���V<$�äTop{�G���]њ���rp	�������I1���VO���(��bˇ����9�N>�#�k,�w3�6�>&^��p��,�3X��@�;-.m�A��DȚ�$�V��.��PŲkW\��W~�A�庠r�*Q�u��f��Ml�ºE���IV�ʈ�̑Vj���0�3���!��l;S'�ZMS�R���j�OfhV'#���<��}�\�l��m���oC�l�����r�D����+��-%���u�o�~�ݨ���~�Km��ş���=+���>�S�7�b��7��������Nt�[�<�ǵ'�+��/<����P����A�2�X���ȹ����V���?��6��,2�U���r@{"�v��/f����#ã�Y vfZ0�#ER��f��`�qk�<���Kq�� �
^��mju�������׿W�VYw�\�e���Q"�o��E���N��4\�Wt���9e>��&�_�I�N��m��V�wz��7ʓ�w<�g��;q����,�IE84�=ux�I=�����Q���8��|Fl��@�Mg5RH(`�Qe|ʶ����1}�'������C�� sKq���)Ɛ�м9���Hبk�ޭ+���2��;��!�@�m���X�)7�X+��#ރ�T+��-���an}��z:�������ig4���VQC/૩
��+��/��Rq`�O�,k
��6��[�OYk�i�d�e#���ꞻ�͒���&�Z�"p-���!̫�l���&��ZM'� $d$���D�N����w�".8q�Q���
��R2�G�!<#�E�A'"+��ǐ��N�٨��%��L�L��f3A�_��NO��?50�/ӑʢ�lm;��LT��]�̷�5�v�Jس�N��Rc,>*B�=��|ʀ�R�/�-,��j�uZnZ_/�J��`_8l󏊻k�Cu�O��UOJ
��H��j��]�����e>k?
Kih��"Ǵ8���ɅV5�i����o��{��n�>��O*��HР R��BS0�������!���߳ ��)������c���C��-���}�鞵�ؐV
�1H?W�䁶L���i��g����0!���!#ǲ6]dJ���z�n�������٣�$O�Alc{��P���f��vG�����uš����d#�P�
5m�w��h���n�U]���a���k��~�3���Z�N�_���=bE�z����x�WO�8/�� ��l]t�@[ ���T��3Kٯ��.S��<e�������JD�x�������48�uO;��!�?K�{��wn~����PMٓ��*�\��Xx�vR$�kYw��x�J�w�&{w�Dw�(+O�A����>�m��;��q1�j�(��{��B�����(���u�b��Fkc��<�Vhj�P%�z�[/���A���ԋ��!�cLw?׉S,0�6o[8�����n͒<�� �~�.*�?`�q	 +(!�����������>ņ"sg�?e��N-�/��<��}�[^��F�P�3��Tz�T����٠���7"�w�N���ӻvǵ'�i#�GJ�H	���_̳����V;���R��^#��4�0��Y�H�b�vv9GohU�?�7Ɛ;��Ɗ�F��N5��ߨ�sP�/j� �ķa����N4W*��X8t�ޱ�x>�I���m-��	Q�J�={F��i? \��Hrb8p���e���P���`K�� k�[� � o ��[� �g��@aG�^�=OΗ6�&�9V�̼(��/Xb��_�D�:���ݳ��B�hu��{��~>ɷ��2�}e*l�W. h<��/@��4�Q���ރ�耂t�j*�n�L+����n�>y�\�W�j���Pzd�cnsC|�>���:���-���p��'҆`��鷏���_�C;Ya����O,���^ �Wff��Y\��D�PSYlHn��V�C"��A���ډg��:-���:���9�k�ٞ��oj*�k9�	D`K��N=����+�����x��x�:������4$.�iL��_��/&Y�U����S�����F�+������t��6����m)����1��>;�,0�UXRRK"���Y�3y��Φ*��È'�q?ל}�%a���,�}�=]-���YV��D�q�)/� �<
�|:&z ++�Vo��<ǣ�-�p~�����捍O����5�W��i��C͟�X��~��赔T�i�N���s��ϟ��b���䖿'b���'p�@A�.;���:���m,@AS6_�/XY^V�8������ox��o����*+G����Y�C����Fs4��߫�O���{|� ��"�zN8j�#�{�P�����j�}�F����	

�ON��F���,������e��͠<c�a�;+�!��_�� ��௷��L�������\��*+�Am)���{�/�'���If檪�����<�H�spp���w07����5���J4�k��F�YY�v��������������:��NVCqaaH�إ9j���(���Ç��]w0hOmy�����ݯ}����H�,//�.�GB|���e��!|���sT��Q 	�	�����L���3���N����   ����h�hKuh�!~@-�"��\ o	�엿�P�;6V��f@EG�FA(�m��es���('�XCK+$��,p�\�AAA�#kDw���^P��X�&gUK$�SQ\A�����ܯÅ���hmƲ�0��?��r�`[W�8gp��37���C7跞)p�����U�����>���γ\{�H޸[Q��v'��oj����o=��wS��&�������=�n-ߔr���"K�~�bٟO�L����;�s�����W+�@X<�i#��9�P?1�N�cP8�*���6��n�� ��/�q[�l�b�_�]�����<�����54���~����,nթV��X�s[Z�V�+aj��T�<W�S��hv�%���Y.�'P��������L{�m��8ׄ��yDm�/9�\��R6a�E­ixh"��5}k�̰sWcB����f���ס	[�t�Ԥ�%7$�4���4E~���9\�"-L�K�h5u �j��9`�F7&��3|���0��v�ױ��Nv��cw-�����q�I��~Rҕ��I�Q8��v{��_^	��x�BR��{��L�$����8+�����0�u��e%��`�Rp����zn�n�@E��eG)1m�������i\�#��(��6��@q�ݥ��;��R�O�Ȩ�l4E	�ye�]4��1V��Ox��E���m��2y�(	S��FS�� ��-v���,�z�ܠ�H��_$��)� p˅�o�����w����	������b��)"	��E��F).!b�y�]��O�u�=�#>G�);�S��5��:�I��c7d��m���_��η4&{h0���w#B��:l����K��<<<��� }�4srr�z\
�ܘ�:8Jp�LBId-l߭�o��>4��\?��K�$y�����8���P����j��t2~�NG>�Q�"��<�����Ԫ����G>�g ����LjFݳ�f�xC
g:Q���1{@�)Y� ��6��,����Ҭ�x	�h�C?lg�7j
�TNE��8M�9���ic>Z%iT�D}O��J	�9��ތ�]����t%�۷^��K@kxt%�>�
^*���2:
��� �PmD
����|^��b'���se�eR���'�Q������0��Y7��]<He�ڶ��%K�L�T��۟9��ok?	.(ѯ��_x_9���h�a~��-/�V�mޱf`���9���Ƥ�xp��@#-���k���4�Ż�ѿSU��!���R�נQ&լ��\�Y���[���b���{���������+/K˧�ۋ�@� ~�{���3� U.ܭ7�qY��e�M��}���#�����Pb���/��պ��5�4=3<�1�^��E�ZyTKD��Y��k�~E���8Vk�\�dg������
�;GR�"�:���`Q�{��*�v+�w�L�N�����DWJ�4iۭ��j�J�)�1��0�j᧥����~z+��N���KD&rЃs/������R�j1�N�{s��K)>8�Z�g�������q�J'�W!�KB����/��UXN>V<����ɸq��P;�:%I9%�i�˪̓0�����r�G�F���7{5Ggt��n��jH�|{�}O������ ��g7k���4TUo&��^p���U���w�����D������3f�S�)���/�������k�B�;����f�<�=����0�y�3���w*�{�vZ%��������>�\��V?+{��5��򇲘��jhzl-�������2�d{�s����y�uޣ��|���'��q���,Ͱ�f��j-�Ct+�RˢU�����a�Oz�$<���R�ec�9x��0偬c S��e��{_�R�?Yb����I��3�I<=Z�n`Ps*����] #���(��u>��E��zS�{��k�����NSLq�텛�_=��zs����w{��-!!q�8����dk��'��|ƶ�f�e]�b+���)�H���:���է�S=""wF�����[߶��?T��j�4�Y��u%f�o�K�^������<��t��q��[���!S�E�J�\�Ͽ�����/�����n���#�R�ae��fV�BEK+H��ԝ����������0;���['���^%B�ʌ�G���>�j�ϊȬL�ACW����n�wE]��t�nѲq�y���/ɕ�"���wŗkh��EЉ|N	�egUp����@�>�ק�>�����w�Q�8��.wETݵ�]-p(3ߎ�t�?�x����%1�ؽ��;,Ȧ�x��f���u���}+���t�9���o�]�JW����ۙY���tt.(��JQ	a"��Gl�%�a��Y�������+ (�Ɗ��T�]��R�C?�9���|�]�Ue���nz����k�Z�9�S"8`�-�8�%�Y�z�����y�B|f{�M����[�M�{Y�y��9��W�e����h�sAfJ��U�Ϻj���D2�}�޽�A&h_�	
���޽{���VQ'��ic�F���_f�э����O��e;��^��#�Qq�9�)*�V�����C��,�����c3^P�/�
׸跻��dO�Д�u���/ɤ�ۚc�=�6U���5ut����U�H̕D!�ּ5b3ۥf��4i���y��k�ќǜK4�7�`�E����P��mP��fpT%�������	qu#[d^������ <�� ���c���!�xz�������:}���~�ue�y�B�c�h�o��
�g�������r:x���ZvN�7�s�E�()�
���b�����s	������[a�"$O�kT,y���{d1W)�)�Ho�d5ɉ�5���8�ZtZ��mf��[|�w�Ia`�"��;ˮ��'R�m����'�7'������6/�����-�e>���O������P�- 
�jrʿ��^K*:A[cQJʼ��D��2.�JU6�M]QJ5eQ�#-Q�e�Dԉ�e�.o5���;r5�!������W�o.���5\���7���y��$��^dq����ʿ/����*$�ɕ4��ҷ`uu�)��m� ��'���+@���.�+d���DO �	]Ee�*�Yi��G�������i!��r��ȝ]O�Ŝ�����Uei�a�a_��D���d��4d�^a?A�#h�b�$$�]XR"}�i��r��ůA�2S�[oO�������Cg��qF�b��
{��m��:2Sζ�ʻW�V|7���{T���ߺ9S]�#L!�9��-^�*S{�>��j�#����0B���Ĵ�=RW�z�����O������dɾ�������O���,'�f`�g��m�U����{i�����\�x����EB�)���9�Ⱥڋ0�w֯���3�Ĳ\�c�f]f���	�OGy�<���Gh�<R�|��_�ȋ��,���47�ĳ D�@�m�{�}����-�C��ؔeZ��a�'6���ڒ����|Y�x��
Ӭ�| g�"s��j�8�������8O�L��ޕ�������i���iH��8�o��E:��W�#�Yd��&��=ʵ�{�15�I������������ª�5��SM����ݻL�-E�� -�{(y5s��%��zC��y��3����b�Ɠ�V�ד/�k���M�Dڴ�i�ǚ!u�WDu��u	�察
��i�t�����ۻJ��(.��=��
��o�H�(R!7KlR��4�p��t{�ɞ���[ݍ�<�Pվ_��em�f����6"�XD~>��k�9@��prp<24d<"|%�BIy�K��
g�I��~B��`��\���~�eE�U<Պ6����3ۯ�c�'t,V�o˒�|��B�~�v/f@��^�1t�rD�����\ĸIx3Q�����e��?~J�'è.ob�r���kʗ�\��Mk�x�b�@��}�G?L���11ީ�z.��MK��S�`���7��k��K?Wz,-�lnA\;Q�:��O�ͺ������IaJ�;!B��׏~=�m��9�r�p!%(��Af�G�Ї�&�W�'���K>�+ڟ�zPJ&��x��溛�#�Ȳh[E�[]��[�7�i�TxIik���[Vk��$�e�A���Q����̣�o�-]�=蚎f�/�W��~��={4�y0by��(5�ğ{?����}�I(��}�_KfY��0����5�
B^ ��c~>IJ���CH����NM���MY7�yۉx�cj��̄A}�Q�_������!�xJk;�u���%I�R���lH#���D�Y�K]8��f��C�|�9��W��e�v�6����9`L�X��L��h������b �]�	R}��o�6z����U��R���Ϻ���yz�"pv	�H�ߠ�485�ٯ��敤��8xxd��%�^�
��#'�[a/��Ǵj&}y�lS;��L.b��0���sJ�l��FImMO���vI�>0�:G _��-%}�G����'mY)G�9.��;��hM�Ic%��&
T�P��m<5��V�D��d�M�+�
��~"�c����{|�w��,-�Î��[]o)Z����)ۇ�$�<��C{���y�,n�� �R���-��*P��/��ԥl�}���^��տ뤪w�����y�m���W� ��v���j�V�����{!�jg��p�2EE�o%zu�2�
�ߖ��й�"�5���3���ƜI��Y��
j��ݷ�|�N�o�U� ��1�p_;] �������L3��S�Y�)){�m�U�B���1���ju���V�)���?;8���~Z�٠���\@ ��d�����܏��.`�ZV��x���\��_:��k�����jh
�����CoH�Ժ����uh(Y'�pc�顡L/!J�)���5v�����cY"�[�4IS��%�^)��6��3PL��ͼ+ۢ��xP��?��׵���z�1�C0wA��lf":����Đ`��9�QW����S�R��e��9��ش�"�L]P��4�-u��\w�#� L�2��T��$�k}��X���i�Q��9�x�����/�g�-/��wtv>�b�I�#�FcD��B���דfwf��vQa�NS���"������c�=��-�f�
��bX��� 5XP3�	S������w�Λt1U��M6{��NtHH���d�z��8(N]����/p��Z-�.?̇\kT��2,s%#0�i���z���l����N��u�+W(]�ZV羸U'���1S�w��R����xa��]�ОX9b�(L	xz�3-�Z�:���=��u��3v�E�P�^i�|t˥g��>��K_�8>����#����=]|���\��36#������9�����;N�O��X'��,���c��&Ů�	#_�(��;~�A���p�Ж5}���~��1	t<����2!���V��%X%Z�bm�GlIn���b�����ȳ�?N�X�-��k��Sqñ�ۤ����*��:٤�b�Μ%��g�!���B��9o��Q��lR�I����v&����#�0�������΢ϋT��(
����]�'���W�c��� #s3���gq�7�uq�(����wUM�=��'�E��`)���������긨���A�CJ�F%��TJ��;��2�P:F��C���;������?8�}�^뉵�>���\r�z9�g���f���0������,�KU1M�X{^|�k\������~�AL;dTHgb�����/�-1�N+�~�D���R�F��xK�};��ײ�ʰ-3$<��NL�rz~~U4��_3�Kwމ��}~RC���7�w� ��?����k|,�E���	TR��pf��r �K�}EF��wQ-*���F)��lug��K�܍�Yat�
�8�LL��]>�� ���G,�x���߂�Z@�<�4�9��W���]����8�Q��0��I�����U�h�z�؉7`����\=N����M�5Ȳ�]rh��d���PYT]8q qp�:u"���>��N���}3b�|�S����u'giG�&I��Z��}ȵ\��b������C�:���r�����6s�؁'Y�bA�i �6	�Z��W��<���fo.;L89�ޗg�?�yS�b"O�0����'^[WWn�E���j�EB�F�����	~rjhxE �s*rb��2�$k|.��{����b@ԙ�r���ҧ}��`�i��xG�&��#_Q�x������|�B<��Lg՟�Z�����	��8����(����M�)��!�Q��ch�z��:7M�ýp3j<���x��T�����W���+7���j"��f�W��m�W�\7��m7t�����w��Q�k�$�v�7��xY�HA�tW�˨Ev��HCu�[!���#���!��~�+��eE���W�=�j���Q՘+<�9v��9�� $?�N�v)����$���A�����ŷ�&�jq���N�s�^���t�Ղ�z`u�Rp��?�=��S��qU!��{Sj��e�V�k�A�j����#{`��_7�r�هA��ά�l�x&R�7 Х��U���H�pOC����X��t�E��ן_�����F�Z���/���yыɟ�3E�=�����g��������D���rȍ�N�p�}+�3�@�qNif�Ә��k����*��v�"�#�d�!À�+k��@9%��¢����G��� �nǎ��K�%]OҒhܰ]v�ClLI��9�UǪNPd*�!�	f`xo����)��j�ow)�}�0Z������������`�G�DZ_|&���69�`ܖ�c���oԏ����׮� x�ʤ`�����@A��ϱ54�����R��%G#��­�S�FE�A�����'J���b-�a8ڸ����Y@Ff�)ī�{4�.y��|��"iŹR�c��Jm覈�N���ؒ��s W����I9NH�e���=��SW�r`s��?�$�'�Irer.�,��_����IiiQ���ii�i?�p�l�������X���W��!X%o��D��["e2�	e*$��K���w��G��I��e�t��z	BV� -�j[��#*�$��uZ_����0���ݕ�gë5R8�(�UL��j�(�?�I�9�Su?uf_�@6(LT}�����E��op��b�e`���2��q�E�ޱE<@M�5����� �k�|?@��8���<J��ȁI"���D6g`����\&}�W^1���X�&�Wy?��j��I�z��H�����9�T|�y�y<�wVd����Mp�dT��=�!f߬똨
j׈����]������[n�G9�ͣJm�lr@��A)a0�e�Nu��H@���LV����/F)N
�
����բ�8��׾:$��!E,�����Jז�ƺIݯH�����閄�I}�⦷ �t%]���n�dj�%�&���=!�n^9Zʉ���P&��g}�|-K�[�@��+��I�=?l�V�1(g����c`/1�L��󽘰�w�"��WM��1���[DkJ%�$��g
a/P�6�do����b�u�>5�a��*����~T��a�ogs�y�ʖӤ\�@JN�t㐂v�+��ʤ�h���A`�[4�9�M���đY��]�!)����P֠��aϱ�T�4��G��U "���~z�_�`j��@m=����]z��c��;��ǂ�n������)���hh�72��Ѕ< Eы�	�4�{	i��x��$��+����V��*r��K߾�-�'#9�Ÿ�?	������H4����DQ�5���mf5�~�tݶ'n�XiF��N�6�����lR�)I[Z��]���������!*���~W@i�@ �]Pڇ)�'I-�1:Óh��WEK�.i�WZI�>#?�!�"7#x�
l5U?�J�i빬j��2X�{ȟ	���i�N��>���T�a�@
��֓��1��C�T�ꈦ��nZ�y��p�Wt�����C�:�YYh��x���X��$h�d&{�Nqw
�RtZn�|��Mv�UvC�n�"��H�'y��������@S�uJ&�N�[-t_�x"���"S�.U(�݂?-���W)�mn�����������k��s��N������44�`��Gb�L
(M���I�u�'����7�����cn��fD�zVM�"1q�[d��9*�o�dA}T����B������p�nu
�d�*λ�ºո�M��1X�����!��A?���W�kb�&�``Jɝ�M�ZO2Y��'����[j��]���>]�m?Lz.��&N�*j����Un?+�]�Y�BD��?���O��X�u����2�ֵ3ړ����}��ʔ<�����`P��q�q?M���)"�G>���9�}��$L����(��Rz������7?Yp��cp��C��`�J�`'*K��&|���|9�Wd���ٽ��{���]�C܊�Q(�e�ζ'�M~0������:ܐ7��IL^^�\S�����8�Z�Q��F}����i)�p��qkLfe{�g!��sf�tA�D#�g�z<��#���b�u�6�4��%%����� '�c�ꍠa�}�@{��^�D1G,��H0��a(	�Ltr!�s�z��*��"$�c8��I�'&<�H���iC�iC�������f��g��j��\l-��YiC_l�=P�FSt�P��f���	��f�!�\o�����ˑ�p���B�w����bl&��VT���\6�\�����_3O6(ZM���K~��+-�P�C��g�|itK���^��z���Mw0ڼ4��O]�O����Ǔ��� |�Њ��E�I+���9�����eZ�W�­���V��琏�T3tќP2�Z�;o?�����5�D|��̀��#��Z�\�pp�0�"`�H@����RP�������W�����e �jz�$��!Dt��X��e������������>��:n. =Yax��� �����n~�P7=,����p̄oU����� �?�#v�?����x�S�K��ǌ�O���{�P���W��|哺&VO��:{"�s5i_��^8����s}�H)i�p��1��Ƅ���n�1��^��������ff�O��%�� Ҙ_��)���V���Mzv.�Yh��,���}j	
�Nͼ$��)��^�qM�Ɯq��<��-���*>HbV
�^A���잻�D�b)�I�8�! i�X������s�,��h��}ʸ:��`�b��W�n��>`�λ�x�8F}0ܫ��Gy[Y��Fs9y�-6�d��@��t7I"lDB�0k�
���E�Y��;[�&�3�m���/�0������=LǱ󢹚S
O��C�'UE<َe>��F���UVr� !��t��wT�l�-�X�1��sd��Ao�MG�X!��r;��le�&�3]����-��&:9c�jD���Yfi�U��B�r�%����o��K���^Hym/࿖��� 5yZ����L<�Mt�h:f�xh�U����>�ӣ��]���Gz2����8���;T:�j>����Z��ޫ���

n8�gffTc�g�M r�9`j�/5�*�;g��,�^������%�n��#ב���Yg�4�f�]���\@��}������w����F��9d��ĉ
q�����B��ɤ6/2O�@:�U?���I�4in}��0P^�S�����/��/��G��Y��+��~��ZΥN�A�X�Q�˦��]*@�s�o-��וNYqd�sAE~Rh6��i͚�HO6z=K��p�d����v�(�US���2qܷ����Mw�a��O��g��j �/p�4H�7��d�Q���r�l��Zo�_�'��v3� ��m�@�4x�"b����j��<6qr"r��~�U��PGZ8[�N��4a��P �� �Y�#�� �n�֮��Zg�����|>�~��q�7z2�d(��EĆ�+c�{�ړ5=�'�Q�9�3I�w����-Tb�=!�x��ĸ����s��w��-hmܤԇO�~a�Ff�&6-�D�(��"�t�m�wc/�2jj���^6���y�G�dq�po�+
 j~�q��T6F�=�(āÞ�!�g8�O6����I��c��_�0�L�Lz�X�˲J�[�e���2\M���aք����Өyt6�6�Ǥ�[i��c8�j�(0��x�@~6�M�2�}Q����hJ�ƺA�xĊU����@l�θ1���g_sG�UMaPq��s��v�S��G� +�]�/o�6w-��/�l�|߲?CJ�4�}w*����n�C=Oy����eZ]_0呐�;c�Vz!d	B��Xfn���3RyY� ؗ��a�/��{֜�fu�%�F,���Ђl�I���;3��	��~��������М$0���W�Y@�sB���rcst)}X���W0�����s,ʯ�䤄��# 8�
�����췳�J^�7�2X���!V��Y�mͶ�v���X;: Y�����a�떵P>����<{{��e:"ޯ�'~�
�	I��K����zڳ+T[<]y��r�G�5���D^:F�t�40	�0k���'WK.���)��;L_�J��=K`Qz �J��ڃ��
����xA5��r�Skv1�����bԇ?�v��IW̄�*eq�����tw�b}Y��S�o �_���]?��}g���@H����{��A`B�	�}�S���L�K���
�"�����{�����R=Yr����ԡWoP)�Q����/�Z��.�ݲx���HB�%
�@��؍%E��ӄͷ�.Jc �����X�|�vy���w�r�a��c8����y�&~/��l�7u'�S]*�%_���MrK���p�r�zLe&z�Dׯ'���Y��=.))���j錦6��A�� $	8��;�!`����=��v�`}j��J�|��q_Dla�r����s��P�Px�ڸ��#�s�e�:�{%#�	y
�mnd��GYD�Dhm_{ٞ�9���<0k�J��M�)j�M��`�\�����e��HA}�'
��ĺ�2xhN4W=���C�H��@�����Ty?,o=-�h�����+�vY�����-�8���ҊT
���Y��G�����Dj�/����?��őI\�g����?���&���ؗ���X�/�vP��u2����*�;&�xx#�� ��c�S,i�R���-�o^�n[CY% U�S����WYm�=o5��
���-�Ơ�B���3<ե��ԝr�Hf���������*n��M�1nv�*c�K_ˌ`�~jީ�#Eޡ�4�ƽy�����t�C̥�c���5�L��z�C�;l�7v)�n��&�վ�_�w� ��(O�0P��P�h@�0B�o#��*9-8��1�F��
��l�ʘ�5m��un��Fϯ� �,��K� ~l�C��[�?[VxL��n��q/,����x���~���!��4����aW�:�Ô�v�����X�� `a���-*��Uo�? 4H��Tr~m�h��v&>ea�b�-��3�fF�F����Z�XV�2O�F�Q����,<> L��	�o@�&�'/��6��S��a��Ao�>��6O���oH��І�W��o:β�x:>��Q�>�
d�4�d�!$6'����䏌�G+��K�h�?\}Ǘ�i���PU�H.۵�����>;/z,�|�	�V#
��=��M��a(B�q?u��((��Z>ʫ����/�3?%��,+{�T��9�1�q�.@��{aa�����@�2�"��uCY_Ai@j�������=��z�!<��4l#/T$��}�^�k�ͣ:W.ÇJjo?G��b�=Z�>���/=nWv>(�p�e��R"�#��O��\i�E��*d���5M�q~��0�����o��̪}O����MTQ�w�t�L2ϛ���Ƴ�]DٲR��H*u�U���D�Kl��P'���+���鎔L�N2 ��Q�_���I��%~�=��L3���--4��9���GAA0�?O ����t5�k;��G�qTK��^�k����b>Sܥ� ���2s�e_��Gw[qrr��oO9��I|6���P#��B��!���{cc��h��"��o�^L�!�1�x�6��P�r-�nʭ��/�^Rs��`0��.=8@빴((�~\��IVE�\�ͳ�/���eƸ�^<�n*3��ڏ/
޹64H���d#�"Sw���w��p}`=�^v4c��/lohWRP2E��W`�T^�c��D�?�`�.���]�=�g��48f�����S༂td*�|;�!�s�ykp���M���=�[��"F)�l����"��8�@��*�i�u67��5�t�.�}���8$DK���#kv1�	b����GKB��~�mg���&��A��csF~*	@,cOj���L �?��Tʡa�+Vz(h���o����r���Aj�����>��M����R�_��^E͑[Jy!N	*;Jd���	�`+� ������3�_�w��ޑ��eH���hc�� 	���Gi9�&b���WN/�j}��Z�����SJJd��u��#��ih�/
�5���o�\s�)��]��7O�Qx�l�>��{�>y��hn�@��؂��?����w!N�~+��F	0��d��<Q~x��n/�  �Il��
'�6,t#���O��HQiF��yA���p����T��SC�����P1�M3��cG���V2�q����/�w�FffzQ�:��ӭ1�x���[IJL���H��A�ݠ�̴�Pt��x)�x�9���E;�_�����#ޑ�^�; �$�!� ]�f�1����{nM�♊�#pQ�P�Z�3�o�Ҕɘu'�a��[�X�B�qǟ���v�~��B�T#��E=E�i�:��� �/`�|_�#���6�>�����(1_c�F 6���2c��vؼ`nnO�p��&��r��\X!`�޾���C�hϠ� �\���l�^�GIt�|.66p�;�x+鳕�:V��ĕj�	�b���9o����ﰠ��޸
0/�k���U�0Y%粦m��dT��Q���N>��;�J�ME�+�}���ո�S�/ՂJI�h{�������t�����J�x��G؆On�����ҟ��\Y�}���/��NvZY���cTv!GrJ���|tY�5.E$F|��)q��{���o�p$�C��	��Ce��̻W�;t)���D��1��ґ:>߄W̖����٭��I^��U���!�_����D�d��.�]U��Za�5� ���H�l4Тk� ��/���4N�tA����U^G�h���D�_�T��,��(��;�3��O�1�"Re��H�nn�����a��:�TY������=�_��z0��YT~C��<�8~OFN�w?�s�� ��}.�b_��]�hǃ����5��ZD<��!�l���WUx+�t�Hp��D�̌[�#<��L�5�����>X��WJ.d<�[� ?���TÆ4Ṃ3f��^؅}�B��F�t�[o�ܾ��:aQ�)>Ⱦ̜�Nyſ/4�A��q4g��,f�P�ł�# IL˿�.�<33��w�hKۅ�/�(HJ�l���$��͇�8o/:���S4�`'*}�sWlY�!!�����o*�z΄IO
��-L�U���kBQ���Rۦ�� %U\��U�������J����q�_�����A��0��"���tdc_�=	5l�	<��Pa�h���Ât�b8��>�/�2z���9XM����e����Q���v��M���L.d�@=����4`�⮮}iG/E�5����-S�/�� ��h��W�v���H�\ �)a_�9�7<W4
83���;:�]���P޿A� f��ޙ���`N�瀩�lo� �����[�lPb��$���-�����!qbbZ$�ߔ �{�v�,I��#& ��#e��d .��]m���FȄ����z������/1�G
@d4��3 �(�D5}wq�SE����PJ`DG}� ܼAl�`G��/����!Nv��pynv~��ذ�}���gn�Sl2?-oO�YAgO��PP��c�z1��Y���N��A�~˯C_���&�?=1rh?��"�H����]���v�FOM�L�\���_�~5o��E��=����̢�!��My4 P��ֱ�$��3݈�B��"��O6�<jڧ;0ѣLv���9�qC����+ki��I,U�~�ϡ�6U�ܗ5����Exݵ���V��]?U0J@5��d��;J=��:���k/��M�<`?*Cd�,�k�$0z>�b�D��]*k⽃�" d8)�!���!�C5X��<'V�����n�,��f�BQ���0�~�����H���=uAzJвnXzŴ|�c��p*�)>�_��.׾�Che�r�v���Tl�kx�<� ��f�s/�Ũ�3C�ݾ��ւE�+gt8{A�R�h�*It(i���$�1}��xm@ʇ����V,����>�.@eL"O\���F�s�8!>��ϜzDѲG�Ee �T�S�������^���wo�d���=?DF�})i=����J�y��N{�������u�_������V؝#�iC*���B���Kvq������.lǨ/x�_7@Vg�j��tP��s��p�/_����M��О�܍G�K���1��ė
��5�� �J�'Z���?ܽ�4�׽G�lx���A%)ˏ��U��H�9���W�G�.rh���9��>�9�� 8�ǡ���b�Ε�D���c[
Hvܛ�.��%�U�����{<^:o0�����y1�����W��	�>����ͼ���6�-l��5����;6��6�U�D@7r�X4�ڪi��M�
CV ����?s�ܖZ�qFܻ���d���`#�(��Ξ^Y �~�#�@�q�#��X*R�AǞ1�D�^Ķα�eP���@�cf&�Q�D���.V��`�;�E������'~�b��ܗm�����'�o�^��I��yx�*���Ȕ���=�ѳ�}����Q'����j۳gP&��\�,?TC���V�RL���+@�d���-�\�_u��T���*S�w�6�it���Y�~d�^�?g�5����}��o�ɼ�p^�rm������;P�f| ��0���i�D���qr�m|���?�1�;	ĻRMÙ��3���XU�s���J�������Q�ß���ˡΨ�1��H�����1�5��a�jN��F)���7�,5GJD�k�d����
  �a�t��V��.��CS�zrb��X�~d[�3
 .��<T�(

#J�jL���ۨ�ԕ�04��G��w� سl�qzIS�w�٠�r�S���	��M�
}������R�{3�hf��[:���������h�^��������0B��̒7]�}Z�bM-�K���l�9�#��G�O�%�Mm��]�_$n��1��.���:f����:kj>���{U��\�vmg�I�U�ؑZ���ğ�<�6 ��k���DOk�#(�;F�] 	�:����Z�9kK(��c3-��|@��5=��i�Wm]� p�V:�?�?�����f�G~>6�E��]e6����B\�)���b��\�Q��k���t��X�k��'�	��� n��&�&~2u(O�+9���&�qQ�����g�kJ~|�s
��2�VLf�ש�֒�ƥ�����Y�?S��B��G���F-#��X;��~7O�T�7�d)�����[���o��C���
!ɱXv�љ�!I�J�a�񵄀�L�Э�;&�	�"Jw�g\���b������I�ܴ���vX��Kg�&U�̇,�{Q�lN�Ԍ�X��{�=�kx8O4�d�/$%Z}���4�a+���]���|@:D��<� e������z���:�2�=!��S�co��|&SO�+�
����XUmrhSu�����.A�6FDhA�A���"e1�OgwZ_"
�3p�\d��|�_�/�8*��_���J݋�2K�%{a���8��v�u�[��`&�/E����\���;u`�e�r(�\�-�(����op�l�{x˪���O��q�,�����x�*[���_��������C�:��()P�^����~�h �>	
��C*�)k,��Z8�l+C����ijIk���k�=@��K�ay�C =P�=nX��2vc����,��@X&u^j�r����"���G�x=���>F�,s�&�����RAC��U�Y����B�%�{��P�D�q#X��g��SN=����u��8q������������y�\Ũ�W�e��U��'��o	@�ii�:���xD:k��[	�<�#��}h�Wx+�-�=?�v�L����(���3�� �hI`��D���?s�F�u������k���{ܔRa���$,�t�}�K�k���ʱ�$A@�V��D��� ����q�.�|jJs-}�����M�K狡���2uO�ߓl�FT) �Qr�6�\��v��� f�C���!���˩%�0��`rKd�I�;���e�����)�,�u#k�q6���w.ϸ(�dp�wR<�v�s� X"���#��Г��� �4�HR?$�[HH
ֲ�*��o.,*I�eV6KO��t��.���ELdU{@�2�i�.$�ԝ��B���t�����=��˨}Vz&u�1�J�Kª~��w8<�E� ���w����E5
1-��E,�bt�OY���۴�lAV`L1�G��X�֏{c��P}�5�hՊXOZ_s��Kql��
�5`s4�9��&���_�j����)��ȃ:�Y�꽪��R� G��G���L��'���Ş]��=N�:�}~�%g��%9=҅�96.s.�E��8��i�E�[�Z����?���7�5���g	c كȡ� ��䀿;�%�S��gR��y;��!��WOY��:�7����\o+NY�����LU���ݫ�_�&���[���c���������N6��TY`�3����
HL8���P��{t,�-��w�-�/����~~N�YO�T�j},eϹ�s��,̋�]�}��7���;���]���P�m�s'H�{#�����1�?bEz�xCrp�ܰ�d=~D�qc�UW��=*�*�s5��/T����m\�x?C��/�a�f���d;��N �x����.	u�n &�DIm�wCɪ�F߸("M�r����~��!�����:��
G-D1�I�r�4�xJ�OH�2�Q�b��ț��[��=q�
$@��^�' av�o��L�+Lw��=��;ob�	#e*"7�����P���]-�*����?�(��2�ÛH��B��X-]}��&dt��$� ���a9$�w����Q���-��`�����H4��~��X;�fߕ���Ͷ�"^kR���m��o'U�%��W�Y�RЛ9�}�:�3ts���mbI��J��N��,���⇉]*>�q_��x�G�3�����̻=�<�f�gÉ�G3����_ �'�E|�ך̜oL�� Xĭ�zE3[.���E0��F��S�ʉ_�	PCX�*�D�\������y�6����)�c�2xKK�ZW�����?��D�����g�g"��G�o�,6��d����.(���:�Dv���z����Q�1n�N��|�¥�p ƌ��]�ݫ��h-�z���wɳm��>[W�w����,��#~=��p�L�sO���9��&Ou-�v�"�_m����MO�+Bz:-�P� 3}Y�t���Fy֝3Ӂd��
s<&���䐲��p�%���=�W��m�1c��LQ�R3�I ��F�\��G�@þS_#Q��Tx ��_DY��`�ϣ�ܯ3�\K����rp��w��ڡ�A��f�B��"��C��NI�����'U�ETӘ�Bȱe-?��Xe\�h����_	�Ӂ��\B�7���a'���T�JFT_�^\��T�/�LK�yJ��k+d����׿�b��w�/�y��Hۦ�-�zh;��%���˽I�0a�β�Zbn����h���O0v��PO�Ǵ�(d���,� �#�,�=&�օgZnUZ7�&#O%0��vHd%|��y�"mC|h<���������l��L��y�-���\���aIr~���$ �6��<���}�f��=���g�Ge&�?&:��:�2Gd�$ �O����.�]��3��U���#ZǢ��K��/N��u�������Yȭز�7���Xb{B��^ƣL9��Y����S��$Pi���ا��� P������{-*����Y�>��6���A�P�x��b�5�u��Z�%A-Kۉ�hSb���&7d�s�.Cz��&E�3s��c{FU�Љ��ӜR����ʅ�嘮^��)��=�C�7���M�p��!��@�B�3�e�S$��������j�z~�뒋&���w�Og��rLty���@�/������0�|��]�d�F_"�@ Քή.~~�##j�w�c��U����W;.����g��t�#I�����H����]a���m���5ɷ�j]�%���r���Xي�aݱ릚*K�y��4=�gT�QZ�z����CQ}@���FA��5��7L
x�M��,Ӌ�}��
��y9�oM�͊[W1�M��Xt J��z�Mb�D�Нb��w�|��+�����[ZM</&��9��K[�ﬕi�k�3�@�<ϟ�������t{�v�� 8ޙ&�&��'.X�E���X�..�,\�������C�RF
���.���JT�����_K��Efa�vn��]�Y&	�<�TP��*��o�2�䚲[ۧ
�4ez2����׎���c��-9ju��.Ksr�n��	��O�X~ֿ�]���5���Q\�_Z<)��C��M�5׎>�������T���\PpMҽ>�, �����n����= �{&�3ms��i���ީ�����P�1>�Y����=�Y3Wa:;7��j�
& � 9��۽��@��0�7e��|�-ߥ4!��z܄�˥G��%&��k]���6Ƈf��9�-ebK㖶D~i�.&��</��.�b�1Eag��^�<����&i=W]���)�z��SC��F*L��9V�CQ��5e��3��^^l�����CB��b2���A��q��Y���hť�3Z3���$Ҋ��EӔm��TKw��G�U[_���h�?< E����OMT�=a�{�ލ4e���Φ�����*��79~'�ɾ�u�uw�"gZ~��g�kVS��y~����J�	�i½�9g�l%�-�]6_��#���24��-&*M�*�~��vrۮ{!�kv�(�V'�t
j�&f	���T�����Jƺ(��20��1_";e#��<��ӶL�̎�$����pՑ�R5���	�˂D���,v�4��Y+eoD�%�?]}�����{�z�<�%n�@��6��_YY��O��6��9�]��He�������f����������~[��_�J�	F�e��ʂ�����u@�{�3�J�T�M<��c����
������.���ELQŎ�W'��F��E�➃���E�ye����ޓ#����ː4k���?��!�>�Cv��.xk�����(k�O�=�7'E��
��8:��mV���0���,��ty.�TX�������ڰ��.Ὧ�z�V3������1�axU%	&�ጴ;:�I��+�q���dv���,���x⃪z��;�xFT���8 JT������ǞQs*�/��q���bh��;��r��k7-hЄ*�}w*
Q�Y�i���\�<�.���{�nk	�G�D�a��y��7��g!Ce��'�׍�2������J`�;,�}�P��.Z�=�����gz�#$P��o�;��^�;z?Ú"�ȉ�����8��j����㘥��,ˋ��{�O��𬋛�n�|����I�w��1K1�����,�{��4�ǧ/)Ws��7��[%����H6��{~�H����6��y�~�$�-%�l+녧�*�j�y�����uܻA6&��<Έn ��Nr~Ì��f��};����-�P��s2�04�0N�V���#e�6��G�ͺ��T�R��@��%5������4� �����$����!ͫ�����	���^7�-֖�������x� Dns�,�Q���[�HF��
_>/X���wR[�,e����t�S�ە)[!���j���<����,v*�8x�?�S^����m��]dRz<�0��-M�xV���}9,7q�~���� �X�!"��y�i��!�[^��'R�KT�N�	��r��%Z��TIyM��7~����e�ۛ���>n��+��5�p������2	a�����-�wN7��x�c��N�J.�|r�>)`M�ů���~i#U�Ej�Xׁ�󹂦�^����<i���E�o8`�2��S��d��O10�r�5��)��2æZo+��DŞ4T�w=��2J��Z��qh"���lJ�6����`�U2��q�Z�nT�ө����-���(O����~�ѧ�u���U�JaM�V�F��]=F��F��8��(7���3��g�K���̴;ߦ�.����L{d�'�R՜k��߹�ۿ���:��ƺ��_/ݤP�~t`�B��ǉ��tغ�9q�[h>yg�����z��L�`�ۿ���xo�~��)��tn�A����~�)a��ӕ��	wC��ߕQ�ǆj3�g��g������rԻ��/�4R���]rG[�{'��`�o�V��w魮��P��}����e���ϳ�*�\�oORW[G/��c?B4_e���]��;����rO+�Y*����DU��O���i���v8��<�\{�w�oFԚ�]����KƪQ(��p�6�@��fi��բ�gR{;�˥ Ih�������wu�������&A�bw[*E?~Ȕ��:�,�����l�ٛ��)7�oc�ﳨ����v*�8a��)�9aI%���?>�(qv?�|[Ԃfάk�aJ�[����~�cN�.�p��j��۫g�N?d.�a��B�*kYL�n6�9�(j5���_(�*MJ�� @w�i����,��Z�C��G��	��H�N�#Dab�g?J�,⯱�������n��ߎ��kԬ�Vq�����y~��U]<�8��qh�m�CQ M�3/(FG/�"�E�����C���޾j��`^���n��.��Eo#�	Zs�����~݁!q%.sG�+�; ��|S��������)��������L/SȒ�zF5{\��{(�i$5sT����ϰ ���F�K�_�t�����y󅦁�b	ϛY�{?��:{Rk�Pl�
x$�P���Pԣ^q۪2($K��d�]���H�"KBrr�Y�(������g�M�h|����&��N?m�����r��Q$���,<t ��dri��j�2H=P�\.���p�F�C��QLa3�*�q�����d��h +�3��^�y�r1l_��V{<�{X�����_�e����b7D�i���J��-�ꎌ_Zyف_�����Ny�"�u�8#J���T�����P���A��m�[��At�i6� 5����hV�>+_��d��TV�ta�3��l�
w�i<;���7В���v�@�lP�ca![������Pԭ�UY���G�9�zF�~�6��w����MCS&�̢ÖC�v��-�
�q��_���a�c���;$u2YP- OA��q^)Y�a���~��/�$F�^*�fNW�Թ��yL��`������gy[�7���b�|DJVwĥ��)����j�Q<MuJ5�l�R#�:%�6���˩ʦy��N��� ���~PL��� ���{qr%V�ty�D��N0י���233�i��7�R4����L���vb�I�Ǌ� �Xی4�=Lq��SZi}$c�'Z�9jc�I%̃g&���΁��tM1�v���RwB~-�xWw���]9��$�l��W���1>|m�r�6$z���c�q��!��m������Lԝ���	�s0�Aj;�
���o7�ĕ ԒGj*8ǵ�Y�xN|ʧ�4�P$ A�?�&Q�S��i�GT�5Zנ���r�h`�3�`�Xڱ�;hm�.��B���������j�U�_���?����SG,��vvz�Y�E7�%~�\�W���*�a��x�%
��=�e�E��˦҇6�Ň�ch����w��+�o�k@d��T�(1�!�F��ơ�����eM�}/�x���)ۧ�}ȣ�4�`�3M�U�Qȷ�̼���/0���e���|��bs�G
�Ozc��cʏ)T$䋕u͜qs�}����8[��nb��ܴ	���⾨���ۻ�l�R�=N���gq�R�o��/���'YrRD&�� �@���>y�4��(u�l�Ѕ�t`%�y��P��@�@
��x5�-\�?�:������>��հ׺G~��z;�_��QM}�]c��C�����������H�tK#%�%�)Jw#� - �HIIw��t	�P�C��9���/��}w��r��gf���~��9��xA��q*~�c�;�nVa#����j�M7^ͺf�3�>�|�)-
��}��#�[���9�)����<c�J����R1Y�rT]fr8ȈI��W��(�=��hHIK[j#��HO̤��������á�����ѹ.��_w�3�ԉ�;E��d�5��qw(�h��4z������_�	;�� 1xG��k=�H��']�G{�ښ_��a�;����֥g@��t!�'�s~Z�&�,/%�;ߘ  �y&�gN����V���3.�
����h�B�V�����{8��a ���&���7��
W��e��k��;}����nJ$����d�x]�z�T���߂�|�����t�Uhc]��#����!BLC���5�b�s��:,n7�b�
8��J��K$��U��G��Y���m��o�ϻ�srp��9��C��=,�1nC��W����aþe߹3g����~�h�������ɛl��O�}�[	x�W%y�4�J�D;hƆ�0�Ϗ ��/�v$����$�����9��贁g�4����v���`�������f1��"��#/�L}�Sax��έ�+KK�m�sk��є�"�N#N��5;�v�
s��szgL�^�(�l�В�}�dlde"P�hl��R����'Y���;m����'{׉S�|��@�3�f�]+V"��l��!�`�ި��-��6��؍�։U;�By�Uc �3Ky���<�w��������W6�M��C+g��w�M��o�����#đ8x�P9"��P�W��L�É��+���Z�����o�#����b$�!S�L�Y㤁:��=�y�dO�N�+�jmqmw�r�� ���r���V=3`)�ؤ�3S�e\�X���,k<=�+��
\HMD���^nx��ާ����gO�p��D��h,�?x	�-�O�(ӭ��Fl�<�Ck�e>�Eg_	��e�S,�E>g��D�
*��[����pEy%�JG~�
*�2L%��;ڟ� V�CgFd���l�Z�>�c�&��-�T����8�T�$;�(иs��Q���7KK�[��h�M�{�
�hl��!z/��.���2��Vtfn��IC( 3�,͛������O^��n$�c6�� *6���������U��k��r�#rک>J�]�>�����b%�yK++0O�x�C�;��S;�6 v��|�J�?H̿o�x>���mi��q<{�;1+<K�"Z������^:-�q;|1+���j�����+����\C�dGQ��Uζ��ӵ�<�ZN>�$��og��"�~ڋ&��Jc�y�g�g���
�L����ʰc�{�7'��-Խ:S�:F�C�%���V�o8.n�5$v7�uZL�3������k�����8�|��733������tW���P�%)(��o���Zʒ�λ��ٌt[m���n�=�ZW��10�&R�Y}�a�jA��Ӹ�0�1y~�N�
�۰o~ ֧1��=����@�!"c���mc����G�.����Kg)���鬮���&A�Xs�R��f�O�s@[�4����wh�_�ȴ�uձf
P�H��(J���z�f�k$(����<8<��Y98� �6�\����c���	C��C���!���i��_�"~�%py��s@�[��G��
�}����8����'�u�O�(
]&��`��h[��+�;��uO ��DD���H.��w�"5=�
P���؜���e:��K�\U0C�.'�F21&ڠ�Jw3lf�ݦ��:e�N�������D8S��;���D�(m��@����xؚ(��\���#s@�͍�DK7���N#^�B���H XA*�ٗ0����%�������� '3�	4������� DX���#��7�W� Z��Y[N�I}/��u<�E	3�Wk���|�Qic�Lx�B,Kt�2N�]����`K�쿹)80D6 Wz��Z����;�����h�Fɴ�Ƿꞔ��LU�E���Ȕ1`���2@�[�����s����vfV�����u�`b>deQx/1�0��P�Qh'�-��,\6��/�텓�LC�j��Y� ��	�yW=�hϗE+��1RRR����s��e�z����%RG m���Y�6"�h��%�w����jq`` ��=����.�]�����1dLҸPaξi�d�<R|#?��C� J}�'%��[S�̺5z����yMؓQ��2��kdf*����M,�[n�w��!h5Ba��,Y�n~���EӬϹ�Ҿ;]g�9g�>`D&d�|l�B����Gd�W"�;V���OSӸޥ[Ih"9�]c���@QFk����W���t����9{N"�=i�q~���/-a���t)���[��� ������V���w�������I䂹��*��'!*������;(��U�Yz[8�'�#j5�K���Oc�ܹs���-C�[������f�}%�a���D{�=qő��L����A��L6�Q�Qb:rcI�#;��Ye�sq�==��7;��ҷc����_�d�:�id�,�1z9�e�9���!������r�K��N�ʐֆ}Q���s��m�OG���!��;l/oo�������� b�rP��=ز��U:5�P_V���� ���Z��$�y��"@*��P�͝�ƀ�f#�v�׀��������˧��GT�+�r��zL׮9W��Jf�ѭ�[��y�	=9�z�EJ�J�g���jz}�E˘؋���O
D��<�*�o*����-����Kl1�w��nNHA^�i����獭#���{�d3�tI�om�
�nYmMU?h ����W찈�:�%H�E��7CԐ�]�@�X���@GC[�Q��Қ���������R����p�>���֑��h�e-��,^t:R���
�%~H�����I1O������zQ������_��{��ť��פ��[�bF�K��:k�|!{0N�yW�� ��_3Ύj��2�U�W�ˍ�ww2P=ަ ƒՍ��Yk����H�هd�k��}]p�QeIDu�R���������$!!IIJ��������ZH��>o$�n�4�ΨaMFH8��$��!��k�㓮�ׁ��9[7���Ҋ"@`��&Pz�r"�=ߨͥGRן4�����M�V_
kk5��X��<}-B�\����K0�`��tO��c��T��a^x�W���]�r0eUF��O6fye���� L:!���Jˇ
0�yW��7�C��UKݗ]�\#����z�6�]aR9��f��C-��q=��2g�Z^vEƗ��<�����~6744��n8ZT��0w�䞞��1;���v�P��ǳx����Aن��������ihm�[��C4�!pf���r��Ƹ���;%����@;[?)�������l�D�gz��e�Z$�� ����d�Jr^!@L��ƛk��˔<�,�5�	���+岦�a^�kѣ� [�1��P�Js��1��"2 �WqR��`��̟�e`��ow$�΂c i22nf�I�~=P���4�2�z�~*(wdo�������&��J��D(�\?|��A��S��jA���{

����A��.�ߓ3��lc��8��������=$TB<6�!����A먶����x���4DGGǘ�NQ="�G5�#�9ZL���@���°�#TTTB��^o\�u���R ��Ϝ5/0Ho��lN�}���v
�4�1춎>��@l�%�7���/��R4/%�ۥFVx-��qN����ùh`_@AA �cI�B�	DP5��U��+C�xg�R�$ײS�¯l
h%�*� �ڐ4�� ��6&���ނK��Gn�����<o	f����qU���=pam\/��e\�/[x-�VĜ_/���� �MO��<�].�q�p6
�Ӈ��9p>vZ��N0" 20�G� ��~�Qw��p;WL�b>H>���_�6=ƪ]�$Ϟ�#��Vh�Aܪ#�%�8<~Kt�,�t7���夤��&0��Jp��}&�x
��P�ܥ�v��f���*��0�F����yˬ׾���ӷ��j A�ٳG��=�!�\ 	�r�:�icIc+��9�~q�t�kp!�3!H O�O��7�}%���?�����6{\�ϕ�mbd�x����2�N��4�`���^�ƣ�y��<�A��A�G���2]ƙq�q*��OX�i`���Q���/e57$����
�7��GGG�j�'���MsU齏��6�ZK1}O:tZ}�?d�
l�D
��r�|��G2$/4O�
��O��#/�2���MMiT2�������0�@42�b�8���r���֮�0���|lb�Qo��ف���nG�V��5��H__;�x��Ӗ��D��O3ė����>�&��T�\�|����t�taB��7N�ԓ���nٱ26�XXX��}<<<�[�v��^�Fؚ����7�m��~9l(����"5�)hg��.�G�Z[�0ܾq���c�p��ȍ�;o�i
�yy�\j��"�~���ҽ���f5����Lz�e��Wz�O[�vD���d�8��~�ꒃ��q

꯱A�d��8��3` #��TٓGݏ���*�B?�d���2w�ϥ��nb����bn���[Pyp����~`��@�ǟ�Q�8�яQd���n''���������<��;����#�BDܲ���uZ?�88rV2|�#�����yy�� bC6��Ah�Q7˄�bE�����9�Lש����|�n���M5U�C�+zxx(�󰡱��r��(��[E����S�?�p��fJ���Gvw?�9�JK��:�z@��I�����;^��٫!���Jd�&-Lman�T\\jn�����êh�)y^s� ��^[���YÅX����zY[���+�yGtӫWZ��œ�R�	\������8~x�
���e�Օ��������/�+Q�Z۱tAO��F6�56�t��I^%�\�Iڃ%y���D��h*i���}�.�e����PSC���:���=dz Q6����*� tK���s>���HR���@M��N;��c`%j:�c���Xnƈ�>����#��z--�I��� �;��*b��2�'�#�R$��-����������x�]�
�1��+��>[��m>�-�߮�9p����h�-�ڭ��,�FW���d྄�&���i�P�b���(�����̻P��7$)6��>c�� ��@=�e��U���� v���,|��ݴ��5��x�šP��[���aK���
��!��^���c�>Jb��CK�
шߔ���H��î7��bM��� ]���ͤR���w��V��s�����:�������+�_/����-���� ����"��=�-d�A���P1��~���Gl�7���6�xg����/�`A���H����ɱ��ފE�H� A�=m�ݰ��Rp�&�UcS_�8���nЖ�n9��au�m�!�k .^�����_J���QVUN�1
.<vh7�o���Es�WYѥ��@y,� �a�E�'9`$)�O[ʀ��ή�[�@O��=�U����^`Ą�8T�uЕ��|uO��ؚk5�k9���V^^TL*'e#��a�5���Apǿ	�Oa��������5!^ޤ��">���t�t�pxo�A��3nV@ՠw�FF�x�%��;�u����Of���11����������2�7�GQ�d�G�C��U������+T��|�+/^����XZX@G/�N�6���	�.�z,'���:��EJ�7����$�z,��BC�A8<?���K3pH�9O�Ș��#	 �T�����Pۼ�VU`֘n��SeR<��ص좏zL�����������2���daz:�21@2Y��a�. pF���ƝsG��&�z߄��<NKC-����?k�^^M���M`J8�<��C_�M}?Z���+D:7�!�<����)ͱ�|C)�G\� Q�ߨa5^m���=M6� 2�c���rr��K	�_�{���;Y[�)ݶt�fYZ����gC	@'[9;4�4�� C�xyy�d�ͅ�Y������j��&B�r�:�%}�A�)��bG���R��/]RR����cL�jgg7�e~cֹ�J"v��J�Jچ�߼��V'H	�Ywi &G
�����'���e���y-���0(��wa�4�%���q��/4�8x��(HlO��7��#P�����s܋H��y��&���b�k�T�{%e�ӵ��M�sw�&��,��Ӕr��ąn]$ ,��ĵ}������R�ٳg�L+��п=F��-����n(@u�������d���]�ѸE�⩇��=�>���2@�Th�x�� ��:I��RF��,�X;���2�n;Pr%���.��wQ�.ll���J#j��)����y
,T��R:�?^��/�4 q s=@����%(Xbs��E"?���V��9Z�Fu�����Y�3��9�ctK/G!(���3��he�𒖖���#��׻tt^��ns���]Vb��T����KD,���ܪnn��C%��J7,��~��I�������2��ƿFio�X�V��oK�L�l&y�����C���g&��xy݇vD������i�l�A�&Z�2~,���� ����P����񳖺�^bku+���_9�VP�|$�-m����>��M�ޯ5㸍�f	��䏛�nF�}�)/@ό�E���$$$�VV�6�4��ٵuff����m��P��m=;;�r��1��,���ЧC)������Ȥ�� C�]�������Jo������&{2��Vxxx�)=,/��8%�IO����k�ptMeL}��f�gK�?Sq#���4�������§y%�hN66����ԣ�>O�꠴��ܳ�ć��s���g�`�lo�܌�pu�����s�<Z�-�V̇P��`��|����weeZ�i��q��g�^���B-S�,L��3i�_����#N\Pb�˖����	(��8��_~����*�,c�6)J���p��� �1�y�gg��3�ffߝ~��������؜:�������22XI�?y��j���ۍ���ө wX=�3�'`�GS�*��!	`���#��&�B��c���)�Ig�N�?(|��|�U&��,�} ��)���w�@߁b��@�X_[JᲒ�����?�*��h���9:��{�uq+�{r���>Q����BzE��������^���\U��@_�����n������{�M���y5j��8�+P�Q������@� �<��g�d1x$P�$���=xP0(��)�B_����VQ*���&
��榚��{]ݱ��Қ��ax��w�;G��"��^hm�ƫ��4u���y8=.�,m,�2_�������*���[Q��w�\��P�����VNBD���� �2Kn��]��_��U��>�F����6�E��p��i�e�EJX���|aikz����Ďì�{2ǃ��W��O�kk�����^�)(( ^Vur�|Q�P����� r��4��7cv��]�4E�?��&h�aL쥏�^3ζ�!�ݛ�m=\���Pu�qY����xJ �*�<V�N��E����HEق��f��$�{��\q+!_����*�*�����(�Rr��g�zJ�#��#�$$͋�:	��K�T�O-hN�9�nn�&^SEw#�ofdy	���
��ڝz�t��nL>X�O�E�i���6S�~���1�i��Nrڨ˹E&Ũ�_� ߀K�j�����a�<��_�6y�[bE-�!��K���*-9򂂗�B�{�τ@�����uK����\27�߷���:�2��PHH�6���S��־����G�������P�=K8���7)�����O�^Q[�ݟpI���k$HЬ�ڲ4��F�8Y>M�A���Q3��K�à���6����K���� ���%�� ����g-{����'��)��-X��3��)�W��߽>9��^�Oo����މM���z��q+<K0�9��7����3�^ٍp�0w�*���{F.��ι������ﾃ��� �/�d�c
h'ܐ̵�����s�S`��5��twx~����0M��c����!he^Fu��P.��G�ed�.� �o��r��Pu(eV$��g���4˵�ʵ�">W0A�cxxg��Qu�_��0sr���;��L�E&�b�?5IFD�-��]x��"rI�e�L�����겇���!�\�T7���HNo��o'�b>�APD��x�'������C
��w����O2M0���O�����b�2��Xߵ� ��F ��� ˈ^�퇍���LR&�[)h"c�p�l�:��5����K��ؗ$^���R�׬4`vh�� �z)"cpZ�{�T�\˺3l���
�(��X,B��o7p���7E,ۀd�e�Gl�X�M�Đ�A\nB��a�d���4����I{S�`C��]���(&kJ�y��-��Jk�����,DQ���Z�--��w���h��H���,Ӄ Rl�ЂG��6�³ #����Ng��axI��Z���N3�n����#	��F�8b����\�p���E:(o.*V��L��t��G�
}��zG���i )�A�W7=�r�0h�H�k`�x�噥"YO_�[ )d�۔n�(��S9"�ɁLhY�fYM���9��<jʔ�>g��/��˦>��'�U�K�d�S�\�8�ʰ~.-%�D���!���\=���[ )���
�����^��>�����v�?�tz��8j�Yv�id4��*oʃ���?����s�[���2xJ�/�P*�����θy�͌�]X���������;ؒ��6%jŘ�p׵Z��|�:�9���=h��'o���������κE�l������TU6.f����^щr=�ˋx�&I	�y	x�fR8/J��{�k�5��Jì�C�#��IVƔ���w��%�bc��
y�K�fӂ��I�[��ٓ�+ʌ�dnQ0��T���� ~n]��y͸f�]b�F��nuuI�e�8K͸>6#��]~jc*���c��92l����﹎w���I��&�ȯ�����n��,�E1��k{F�))� A���K?��,�PJ>��.��Q�����&@U;9��y`������1�gx.�[���ǺR���-]qz���ԁ��ԙ�欪�P��C�N�L�]���]
B޴qAte�T�XҺ��c�CN�t�&����Ƶ0����:������g���ɂ���8�E����T�j�*=�u;�R+9$$HΕ@0��+�HH�IB���Թ֚����@�c�/2�_}O�^�s:${���h(^Bۇ����||N���� �Y�ԯ��Ȝ�I�;��_�%w7잒�}�z8�?�'DE�+_,+j��2%��Q�s���Z�j��-�C�:&��ȱ��.��5J-�in��ʢ�)�'�w����P�X��R�	�}zd�Uզ�5>���+�Vѻ�c�x��;e�˼Lr�G%�,�Aᳬ�ni-���������j珘n����=1>D�{R%�4f�1�5��K�ϳj�v��|RE��Û�lB�tsS�y����j�����W.���/6��cN���Y�GK�E�;f�i�/#B6]����n������v��Q	�ѿ}�"��l}��6��A�P��H��ZJs��H�V_���l$^-��?��X��W��t�|w@�75�nFV��ωԛg|�j�`@Q$��%,&=$l$t�����S�(��u�`4]d�&�'d�G�o����q�?>�
��_TSx��g��:��=�mRp1����^D�U*����_�ñ�oM}����ΆQ6��2�����}� C0�+o�r�}NG��4m=}ve�^R����w�w�v��o}�����i����Y�X�MJ�Y;1P8��EJ���c�jsN�5���eNB�ߌm0|+�ۻ$������8�͓�?�N׻��\� �L�;��0�c���,��(�S��p|�ʜ���5`{DR��2��kԜsвZ�!~p͙t���N����'M���-'?��jrz\���D��6�����Q�����%>�]~nl$ZMM���ڹ�Th��1���p%	"�V=V���=
�,��e��0?����_~ԗ+lp�ʴ�O�O:%���Йoz�C������g��HG��)f?OuĦ4-�X63"�$� h�?!]���^�HM�FQ�m��׈e����/,`��D���KHJR��J�`�	@�]ZR��o����xz����������IvV�i��D�[����s��m�{ٴh��\!ݺ袹s�Cn��Um�sL�����+ � .//_!e�!@��&8�Ü3]w�C�ϣ43��H ����N�KHD���^ZZ�r�e���|��Q�oT���(ŅWI��kX,a&T,���&�W>�9�~�V�|�-�=44.nm�4??���rWBJ�9���5?h˴���֖���(�k��DDD��u�&�𖉡��T���*Nܟ���N�\1�<I����"����q-�r�N��p��5�;�ql2J�[O���UU�����~� 9P�%Y)g�\H�too���D��o����Nd\\\�<��B��;R�t͡�u����}�~I���z�KP|씠d(�aƚ���#$*̒�v��C^%�޴�V�q�]���9CwaI<���Q�W�X��eV77%@l����w����t�����#��8ݟ���L� �o�K^��|I	��m���6"s�>��.!�M����fRhh��R��(���x�Q��;�?n{�����p �Zfyl|<;/�N||��u����j��"�/z�*��}�)��ەr�Ya;�!JF����Y�1�Z�]��iM|�p[T�ٙ3&&�]zz$*>9;�#n�G�A��������������Ȋ
���Ĝ�\��].�^�웟.���Tb5^�a�B˥��F����{��|�Pי��ꇉ�
ntj��P�G�TT�`� KX�ß{xxd�Y"�>I��,��M}ਯ�oEHGG�+��72P�F��(F�.�/3���QZ�aqͲ������J�wd��ۜ�R|�V>���wycccr

�����%��)s�+M��ss�@��>�W~�Q;�E��H�.�e3������r�:�q��ylE�ō#ﰣ3>�A��D��*N�4���{ڄ:�ث�U�RR�===`>��r`ή���{<Zi̙���ܛ��EFb�
�����&=س>�����Tޟ�a��U�`&h�Xr6LI"*�y����Z�s�]���F���Opg�UL��C+�?�N��:��+|�q��$�"alL�<�u�"s?��{Cè��;���hWa��C�����>6���ڊ]��(w}�8��du�7�fV�O|Jg!g���qtt|����iF��Q�:,4TT^�t �I����^���M1] tyyY����Vl�S){���QRl�h��b|iz��Y�t��d�C|���1u�.=9[�Q��{���8,|���}�\4F�")!�|g�9I���)r\w����1����z
ۇr�V)�451-(N�Ho��e�kb%��K���DO�-Ĝ�xLz��׈���SE�����&����5F��j�u=������`"	&���9�f���rr����3��M��M�<��e��o~��>�� ���~�E�w�	s������+vVY��KN~��_���wqᵸ���:��;���q񮬬,��0R���C�|� >�y��r9; |7�Vo��$S$I�LPK�T�5�k-�� v��!���9@/��1�x.HsKK�g��M��jk����,,�2����3̼x�)����ɘ��d��N���m/�,����@�a���rww��Z��R���ۏ���g|�~�6���H�b����� �����[���8|�χq�J�|���S�s	<=����T�Y�dR�((���[ɥ�n��fgf�F򕤍�?<xv'1)��ɰ��7�����
6
*����C�J|���ũ`�k��W1-G�Qz!Yśaˡ�����Ŋ���K�̽���U�g>�������S��Z��_2���m�@�k���	cv��
��Ǡn+�����,.��?����>�mT9����2<İ=��;ra�jkr�wH�DK���ˀ�(���or<6�'^\\ɺ{U��4�Mz:)(ٞK'|i��
�?�����?;XM�id<�3����~����~k;�s�Se��λ���`t44H��$��$;;�)��H!&�\�DI++F(<ZZ!�|���&��{���M���{�bI���~�f�vv�j;�T��G���5�_�C�n]��to���$�l���_⣐��V��1�Z�Wg�����G��ض��U*o���
�����oj�Ѕ.�m�k1g�M�ؖ\hT"w�<ƪ�xr�!"J'B�,{y�8�q>\t�l�Kh������1����Hb��j�s�±u�9�bFe=��55���T�$�W&��e3S�{r�5��a+�����N	>@T�t�Stl�B�s3�h�z��X�﫩��Q�42��t�l=��t�^t��k��I��p�,����}�G_)��(b(�Ia�����+�+�iʞf5�&�� ���+ʅ�?Q�v��سS>>&k��|�~�M�Bmmm�P<�Vv���H�we��L'��~���s�W܊B�?�S�"
|�l�İ4���Ո(x�$���e�aw;m훰��������h̚��'���EH�����>ɗ/�"Ʉ#����\v
��KW��:BR�g�CC����F//��/P�1KOcb��z_�k��)�q���R03�k�9 m����ݲ�˯W.*���3� ��B�+�z4/`C^����}� Gh��Ej����ݓ�i�?,x�����)���D"���£�?B�Ȉ�H)����e)P��|�w�d���J��i�GB�����D���4:&&�Ouk�#saA�d��y]ؼ���(�5A��-W�����宮���p֯��Nb-��zz�� _�]]T@Q:��w��>r�8q�a]�r<�&�������P����`��+)���p��� �4'
o�������r�SG���
ç�|$	,�a4r	�uu�n�_@��8޷�iL3�=%�:j
{S='��N��PHQA�@���6���?i��������'�~��D����~K�fR�ؓ�%&C� K��\�h`���P�l�ԛ����b���P�or�G���	�̬�y�H��U���s�+!�gӾS7�9�J~n����%:::?�0�����܁h��t����G(O�}���hr4���N�q�N+����u9
r�N3���kp^l��^o`?���.K�Uc`s��+֩FED���k�ۀ-�=B{��|l���O�6p�PB+�	���I���=�GEy��<b��x��T��$��^� �!v�Y��iA�ѫCQN�]�n�	?�����6S��I��Y�-�������;ý}�E��Ǳ*��c5Q�Y�߸ێL�V'� =����5�"���`>���Ob�9]��\>�,*Z�ɗO��cm�]�:�kSQW�S^:��Sc�~�>`*�Çے�����G�	��9{�z��Y�BM�Dw��9t=��s�_�!"C��a?�i��D���ZB�k�i���R�}�m�����J�Ԅ��5��[���$0����~G\�e8���0�(1��R�0��쑉K��> n(f��}�=g����CC������-�r��������;,̍Đ"1���?�r�)_�r젓�����~m�׋�Ť�e�	�1H����~�òCRS��S8�uE�u� �{7�m��oT�\I�;!F�Y>�aV��ĝ��`���问�Ej���5{h�b��5��%%�0��@G��(���{}���S:��'~�͎b-,��UL��}�Y��_���n�����?̼��J�!~�!
��DV(�л��\�;|���"��(�����nZZ��i���H�YzYʐ�z�*��'NBt �?�Q���n:�}c�_��~��ƌ9��޾�Ty����Q�y��=��<�o�]�
xhP�O�oC=tϗ�~N����/.�CBC�T>����~߷�X�L$��"zNNN�Q�,N8:B���|o�X_��ج:Ռ�U�^�tP��Jďϱ݊�t��K�R�
������	�ne���x	��R�үY����2Z�lht����� �ɽ�
AHC���*�(0Y+Jo�!u2�0>�_J�a<(�͛5,�	%���.���;ctg>$A�'��UnZ^齆1iOt���Asp��K��q,�`�����T�m�{}j�)̜`L�f���-�=n��n7�.���j�֏��*�����9��
�YrA� ��֣�}��}�����]�8?����c�/��%O��#;�1��k�gt?!�`�EP�k�g$��f$9���h����'S-A�N˷�ẑ����Q���r��3K&''O.�T���ܳ�r�W�V���w?��&��k;H��67������M�Л�o�wo�t�p�NV����i�{NL�`�S�D�fa�s���k���^�,'��v���M��uT��HJ��L��ۙv	�P��𯫜����n!��Bmj$pB�O��鲛�����^��� �UwyWQU���sqq!]�o�;���A���ХCR��%0�Eu�>�^�;�6��HS�H�7���S�e|r�����s� �
JK�n�4���5��������z�����=�o;�,�*C���+��'���>�@�y�E6ѳ�b������^�o�i�{���-YW�˼9{6,��բ���4n�<�	����a�w�P^ٜH���v���w	-spq���g��Rt����x.
����bï�������H�Z��S�f��gcHoƘ�?GNM���r�>!Y�R���]{�.�������d�Q��ɀ����U+��u���oAÔ����1s[�ga�p��;��?)3���(X#�E�Xb�52��r��'T���T*6����v�#ԼΣw+^T�ߑ�o��N)��Y:��r|D�����*䴟�(}4l@����p�$����Y�Le:�$�ņ��_�<�E�$4�t�(���0���X����*ue��K����R���#���W$�V��<����tku������x�-�^H����Cl�\+W�h�ɝ@�G�uk*h���;x��=U��z��+,���-#g���\�J��{{zځ����Y�1^�u�n�+Q��/���߽斖�y�l�6VKOn-�6�}�s�J�	�7�M�����k�wK����Iv+"�������=t���-7at���d�%W�]TԎ����c�_���m̵��ב�o���օy>۽-�[z���֩i�z}\IH�`
���n����#�α5Q��`=�n;X�8�Ǳ���|/,����s���A�r�	ޠ|Z�W�j�1~�!��f�M�vC��5к@��[�1�d���O�WZX�|�����;52�_wH���CS�o�S�5 ����|a!��Hr�w�>�
���u䷕4-�v0l�\���~sNª��O\򧧧I��<����:��8knw��H-o��S��G��wO,i�m"<�>�s�/#+�y��}tz�v�s�/K��{�񲸸���� a�f��lc��ϵ�|���cy��q�F@L�J+��!�(��>����B��P�S���`�̬����%�C9����Ƴg�pϞ
S�d?��u쎇�5�6R�����*������� /qpۍ�- �Xئc�Y��A��e�JјV�+6v��\P��1j����`bv)pϼy�a�s)��Hk�Y{J��R.�k	3�n�`������f�zL�x|\'���&�\� �f�ߠ��-�)�N��A�~�kVC����'I�o.���Ѝ���79E���Lq�ǁ 7�ֱ����_86bGQ�����|o��
��u�w��B����9��JF�����8	\�oD����
Z�F�f｟Y�!���a�L{���e�7�,?HX|����}�B"o��*뢐�Hhϡ���˗`ʃ��Shc�uvvv����e&ddD�}�&p}�O�̼��"g-�h};"߯I��>����!238}B8w���$O�c[��q=�=�Q�2�tJ(��Mȁ�H���V�Һ��1�XDh	@�ORv�?�`"	*�e���+���-�G����#��
�E7X�Ơ���-}x�I:��&�����	^� �ң���]Lȭ48s�L�ߊ@H��p��= �\1��sQ�	��V)�/Q�U�i����BDW���.T�]6�EW��"��~#��4/����k�wy��wZL@�hs<''�u��n-C�20 /����}X�q��)��bf���>*`�r��9s-��_8K�]x��Y}�Y<((�d^X�ؑv���6`��]���4�sK�uZ�L���9��u0�@�EAJ`��w�_�?.�1�����*��[:�s-$R9C��)<{?��5Iw�H~9�Ld�t���u9���܎n����VR�R>Pz�һEo���s_��^wSt�|��pͤU�y����.$2.rrWy4Z��� ������ZQ?��������d��[�v�U��w~Y��ꞷ�ͽo,�f�?ź��'x�����?j���(Qq��bO�G�$��j���3M��yw�~���i-������)�(��,h9�E|�L?���P��zd O�*~��齅�K�.�F8��8t��e�PX'����d�T�)�����gi>�v�/��C��jU[���Π�)�8(�g'����))J��%L��K�
ls>�e�{��4Ү���r��;_:;Oy��W=6�slba=Ɵ��N�W<��@A D3t0T���|�/�%*��9n��C+��}<���uΣm_TX���Ə"��E/��l������C���g��B{l�WύZ�ba����� T]��C����48��Α�eϲ�"wsG1c2�t�?���J�K���Ç�3.��B+�FFFEE�no�e�o
�k�ó�邳KhK��4�'�<*G'&���HV�:,~�M	�7Q�H���	z��}}�ax��j���,���
�-��؇e6;V<�ݖu%$�]�*_�Љ�/'�ϫ8�����g=�W�g�B��X%�fd�Q� 
��������V��k�s�@�k5{p�ZVc�"a䪆��<�z�����HX���д<p|��D��U���_�[�q���=?�
�6JĲv�~�����1�m�� ��\-`�^n]{����z먪��_���8t�N��D���;�	E��� ���%�������{���d8{�91�\k�H��d�6SR�;'ȅ��P�5?���/"�t�+��eRg��]o�g:��Qi���;d((��R}�c՞gf�s��/��F��ӷvv6W�c������ζ�nj��	�]�i��h(�xS�'�	�����z<���"f���rbb�q��㢌���t�A�M)}}��"cc�S����6-��#"m*[�)��/oz,�e Qc"~�O����h�^���Dn"��+ �O<T���100|3X�������
�^���x����EYpa����Rr�l�\A��<���l��j���a,�(�"�t��ܟn�$4,��Ċ**G�0�腋�dߊ�����at�ׯ_�r�᎑{(����a��i+e���ݍwFB�V����]�w��8� ��EԋU^���n�� ���a�O^�qb8u]�����\���'�N�+v�H��mfL|�����n�;s0aO���Z�D;c�k�����d���'��q�j������r�8w�%/���r����P�J1����g߿��O��z�Ժ��'vc�w�@7�qǭu��ohh�a����	����������PI��t��%�������]ZIC?�MQ�9Q�|�}#<����>j������q���� �_n_O�iVW��:�?ߗ%���$\r���|���$%�)��/r��)�`�w��#4�ū,�~��@�)k# �����wm<�hN��y۩���so���䎌�J|h��z_�xq�|�O����H,
x�W�J�����סEC�_���jk\mr���ui�����W�}�.�Հ,dL7@����-z�@hA=������_��_^�,ں��o~0nxF����;���+Qh))�Z'i,^W\ ��R.Z��ԕ%�|"a�KD�� ����I�r��/0Ub�p`&�s�/үa�����U�ݨ�`�h�~��=$id��K��X 8c)�FW5���;�:��T+lll���ݎh��oF�p&#J�)�unl�y;����!.N�����2�q��=WQ �Y9�1��P$O��U���
�������zw���;�ߜ���<�X���� /l��#'ߥF'�j3d��+r����@�J;;;�c.D�+}��Z�Ϝ� ��'��<��,�[J�K4����S����6$څB���r�����y�9��Cw��y��*wQ���4.phZ�}��4��|�j�o�,|�9_h�0Z��fМ0Z5��-��9O�.��M��}P�*��RS��ø�5;����X�>���$�nc��+�~w�4LF��o�B�=�4˦a���!�%�٢�iNwB2�1���(�H�-Y�'�\���r���`��/19����Du�K����.r�?8�Cb(�<ɶ +	 ���p��u��X�W��ͧhK����������|���-)>~PE��i'j��ye��������u��m��|1u��;������i)�׈/�}�x��6���6��Y덏���������*�P��QI{;�L&=��0�ri3��T~42Z��^KIn��.M��/e��9=j�*�C4���ɝ�X���ӵ��f��8��}=�7���2D\��lm/-Q��F� ����߾�HH!��5'e�R���Ӻ�^ڢ��y�kg���rsss]{9� vi�|����-HJx��#t�R��(ȱR���+��KGo����~�ohV�d}�9ө����IJP��llN�[�aS������jj��;�a��:C���عM.l%.R3?���>�u�Y�h .=l���8O��e�Y(&��5�g�~��	%�U����,�o���IͶ�kE�Ԓ�� o�^��"��`0�X'!��[�П,x�*�id����2���܅p��G���ߨJ��!�p�[�hO��}.jv��Ƈ,n;��#<+��f2;1_2�����	�N�pb��(L������}Y�m�f? 1��V��1�n),�w�WH&�98�1��L
�A55�c:/������^��;> �����<v��@�ߗ5{��1�؁�|Ř$jQ�ޠ�D�G��!����3)��
��lQq*Q���G��h�;{��d:�̈�3���3��s5V��z�(��*�TTS�;jX�/�������L�Y�[px6Ľ>��Ո_�A��d�JBW'�@�_�������D����]vE�ϾO�A`�P���������	���a��d��MŴ��*P�yQ��|��)���Eڧs�P�m�K��}�M���n�B��(LL�
����~G(A�3u�F��NN��?=u<��A�!�|s"	1qx�IE��HOOo���]0������>7�ٲ���Ѯuu���*/j���k�Ȯm5Cd}�׹<٪v��tLL��ғ�gֱ�)����T���TWPZZ:�ĺ(�\�:$W�����)#����A�{���:�_�(��)[�#Z����Omzz{�s�*0��9~�� $HW(:AbN���9�3�Ъ/��ぱ�����0�x����\�H��.��b֑[�%�h��*��/��W
aHt�p����5�> �L̛�����Gǹ.QuW��<Q���պ�O$V����q��n��]�JG���ŗ���"��T��A���BF�7����ҡ�"�HOn�\�j	D)�i~�0ڰ��r���9��w��[��t��/V�fN's���Z�zO#?�U���g%���N���� ��
Q��KCӯ��Zw��������S���K�^yo��J�Ԕ��7��"#מ�t&[��!�+�����_[��Tr�r0����0�Z�Q��g����S��0h��0{R��`�����۷�r$R�E4o2��`�F--����-�(q��'K`�2��a���v�n�җ�P%wO������EO�� �zG�lv�;��d��/�x.V���-��Z���RY�p�ka�BT:���KZ��� F�<�%Rs��U�Ȼ���F["Bm�����|���Pv�;� fL�`�NBd^B���Ng�h��ѥ���	qT�¿�
�����p%d*~��W�e�X����ETT���z#�2��y�¶D=Ry:M�i������ܗj�Ҥ�/i��bTf-NO#�� [,�\?��������\�B�4G-���ѐ� ��O#�K�����̃����ZWY�9`� ����e#���A싧
��=�w�ݪ�7�;8��6�a;t�$K�%u)���lؖ�Y4����ǿ)�s�̓�E��[�sttt�qL�x� B��+'���.��S����'f��#s���g�YL�
'q{{ۯ���a(�5��H�Vm犺�q��n�|��^�����rH�b�z��l�u ����,��$e͵��~�]��m}���|���ɇ��x�	䰄ҳ��3t�nn�pm:�6v(P�
�І3�[7���Y�o|�e�����P�+N�� g��A��*�Vu(�b�A��hBZq(����}EH"o�G:tG>m���j��6�� ����I�����w�I %niJ���=f�t4��
d���$$!���d5�GA�n��"�Һ��M/FG��/�V�D7���:�4Ti�VP��^GwW6����F��"��+�c<lU@^�2���%��\�?�gY�4t�qeєg���=���c#@;��沐Ϗu�B�N��Pq�ũ��]�0�3���AߵX�ߗ��[GGU_�<e�������0��`���ޫ.ّ&����ַ)CP|�罴��XF�1�2d�Ǐ���T���,�L��jg<2��)�I%|Æ"�����!$����H��F�H�[��mXf+�h�b�s:�%����x��1@�N���(<8�۾�������U��0@��A�Z�:���
�q�I=�繁�����'��U;��u�)��������<~s�000�ؼ���;�u�����Z����w�ҺX&�YwVu!P}�2kl^��ɕ��6p
�yV��e{��8R��0�v3�
���d�͏��F�ER�Py�R�to6q�8��{��L��;��Yב��ʊ�����*<��~6���5���+�Z��Ax� @��Fv���\\�
	�G.=�!jx5{�h��jLC��S����$[]�����Z~���8����;���ިYe�)���e2�fA@}�Y���3,�_�ˁ �G�V�O:��r�o�v���ػc�fP��X��D�h�6���E�ѯ�tL�E�4S���7�8�E�F*��K��q/�����3J�T��8��H0�Fbe���FvbL���o�����߾�J�����Ǆ�_x�O�t�|(?\0����\N��l�+�tc|;��Zf�,~�΅���zn�cs����8$����/��v�h�X����H��"���9��f| ��8K��.�u�*�K�g�PV������Fb`�}!�a�fKvtry��F	���l���144��di{$�TK}�2�'��=����B��0���6,p�g>��KGk�f`�R'u�X-��x�>}�*H)��~��!�w7i�����O?����=k*�0�� ��d87���h<�܆F@�6+�up�R�v��0�‎:�	�m��o'��f8�qF	��l_y4>�꽂�t���o�F�Uqa�U6#3<����UGͅ�ƿ��������p�)����Փezz��o�c��~����N�OI^�!8��8ݜ������F47c'MrQ��W�{�_�`,9qg���g���V��Q:w1N������W#0�FFF��m����3��F#�G9��*
 ъհ�uXay�L�Y��s���$S����n�dz��O�aSl��	�}�m7f/���' �,�����w�TY����Ĵ�p��k���	�i��LR��n:}i��s�o�D�d�*�{R�c��O֖蚶��M��Q�͎��D���� $�g)G�~�������{�B��o�~��W��Zl3#q$�Ja24�0�Aa�!R�c�<"���S �*�P-��C��Y��b�V�J%����%�Gb�I���S���/�){#jI����}(3l�+���bR301�����;WOV�NJMOg``�^���r����p����C�я�j᜖�y	���UBi����L�W���qs����3)��M�A�s�v��J��� �-��EN}�*��`e�g~�ޣ�Tz^�i&߃k
�;N��޸���O�<cbwOz��i=��$��|�VU�O �*~�=��wǿS,s���{{��/��32HA��$$P2>�g4�� ^ۏ�e�p&?���O����}�nD�2��3B_e��o5�|��X����O=����jg��T'8�t��Kdx���HM���7`�0a��v��7QE;,!�q�هD��dD>T$P�ľD��L�y����m[-��T=6�됿ӛ��_ZQ$9��F�^���NF{a,J��Ą��I.�E5.~�	��&r_��s&{-�4���2|2t=ɖ8��3�Aڌ�9�����@2�5���8��;��_��<�+q?��!)�E�b����藄��=�Y�|���fJؒ.O�@$!X�/�"��vajBT[SUB�<�Ǌ�b�$��2?���Ʌ�U)��X���ܤ-np*Lʒvv���͆��,�!=��S]������.��|�GsVzR�m��3ާq�τ� h�����K[bѩZ�n��f e���!���aB"��Û�x�6R�
��C?��S�]���GW������j�A�$�4֮���jEA��#�F�JW_Q�YyR���9߬�4,D���V�v=M�>�=��|j��ebzZ�+~! �d"pn����ꁷ�Цe���FM�v�/=a�y1QmE��Yxxq漿a`����/|ն�/�) ���%�J����w����:�޽`c� e�r��HV���h�0����4f�_��G���1����0j�{;0%&&�/#���d�x��E�C���S��I}C�����}�#YD�����u��*� V�������i�7�q���-]S���!j�"J�
%��w}P_��<���w|]n��S�q�lB�|y�6�9��$	��7
`Et�!;Z���s:�5;b�Z�:��Q�D�����ӟ���<͓�*a���c��g�������(�h�Li��V�5�w��W��C���$�Vp�C���΄�Z����bc�N��/cj���F%C�	x�|����Y���!n?�)�+w��޸���<���42	l�J�l�AQT��k��0��ܘ�.a ���% �x������M�w�=�#�~ư���k��ڪ|���ƽ[؍qJ���� �O1Lc�T3+�K�u�ؗ:�N]��cD�umC���Xԫ��=C�\A�MD��A�_qЖRD�В�"kv���G���>>��ĩ���%�ޅX���O}�Q� �� 	�i2�n},��:di"�#Vu��dĘ'e���(1����M՜WdGGK��/?�ج�C�19����C2�����m���e	^�n5�>�x�#�$��/��wi�E��0���󋘃��?yl[�dR�[Y%����$����k.ܼ���MC�$0A\;��S�L�t��ưi[)s��M���HWPP�����U�
����KQ@�܂q�� ��l{�}:�k�"��` �����g#�@�ȑ�[]�Sԫu�c�����Œ��>&��}R��'RW)��Y5���b�]�	��C���JV?����"n,��j7��=�\5$1��Dv�&�I^K���M2F��Wv_и]"�	���2SЎ|����Ew�֜���қ�g�$�Ӹ�m�(���s{��R�ECb�/3�x�J�$F���J�����uH�u��|����j���\d��A���Y�r����8Z���J������v-�_��Rh�NPѼͤX�\���ݜm���c)3���c��;���������.ڹ��>揄>�&]٪d���FIuEm|�tL���>j��b�Ng�5��yK޸Z�#f����{���4�(1:�%���8�_����=�5���I;m
��'�P�HڋkZ�v-\�u�!4""a���Uz���:��M��#��~v���J���.6�KKt �C�\�b�H?��Ks#j�(�I�Յ��RNFF����-�Ĝ�Z�q����2�߫ݨ��Wͤ;4�+�������V��~>h7��k�Ң��r�J*6�I���1�Sn��S1�������~+�.Bm��M����S�uJ��׶�N��;����#~�.n�<������~;=��<�x��������n��.��l��c�;���y��HO/Z��UK���/J��oY����i���%�w=���7��cT������{�2�bs��]��E�Έ����@��9]�?z{��@��r����N�OŮ=�9ۂ�>��^'�uB���u^�q������Ԏ+�� �.8�*�$��o�$V���8��ʯ�NO�:�+k�hR�lB�!��~5���=7���w^�
���Qu�×^�;����e`���^`{i��%3l�n���'&�(q�am�A��6k�V$ ��8 %wn;�V�̳�����}|���Z
@�G���u�����ป�_e��x��� ��Z���t��곯�W ^X�|L��P8 0�ǫ�̙8[>_���.��Lj����ȥ�d�@=οa61OH�R��_����r��kbIK�J��;�����/����w�d`o�l"B�[qg~X��Ki.�����0@��o^8<ɫu돗���$>-�g�!LRDjXvϴ+�@	o���FI	�i�y^����xnf>7����t���V�����4z��R:[����D���6X?�!���r�ʢ/�
�ƖB�P�������vY���vP�M���9�������:����h���Q;��|�OO<�sx�dm�	�Ɨ�F�_��t�\�*>��34C�H3�w/ց���o����#�A,�]v�[���#_Y8��-qb���=>��CG�QrJ���м����{���87�w'�+NBxh��2^���l�=E�bO2�'�B�)S��un�(̽e���;��;�*�yZ�}�ϥ#Ę�n��

��O�g��cc;�8��;���Z������|��u�=N�&b��{sZ���6������Iol����Q-E%%
�-f�(�	=��Rz������|���f��=rg'E%F�~/����U��k(�ۑ�����.�&��)���9��<<��W�Y� %��8́��F�<!��%�=z�����F'S�%Jp'��K/�8�KJI��$�0��d?��*���>��S��1���s:�[���A���}��/�w��DE2�*#��Z�2���ʱ��֨�^s���[������Bl�ջ2{�	���%��l�uǂ�%���n:(�tD��������C�w%�N�z��(�ꩩ�jU���`���:p���l�|�=E�~����P�U�\�)9��Y������g0�Q�LNV�q�����W]��J��?'���ݴsS������gf��� ���y��eg�s!��/8�.����꒴6m����������Ӡ<�-�.<�p�	�;����մ6%�ڶ8Rp'm<�X���u^EŨ�$a����a�G�&U�|�C�7�2�/���x�M\�U�����é�4�Rl�On�IX,;q,�zBo,[ք̵�z�?��/��u�҈��������ޠ��^ ����%�ǒ��G���$�|�'�S�l+� �Ó9h~-���sR�?@���,�l�Mx���T2L{��Rc�9�Qy��x]��WV�Uo�H���B���hhi�2*��Z�ir;�!=sGz��RJg�.�O���;�W��l�	����y��=t(>��È�3�»w�&��BB�W����/yoc\��}��r����G��b�������N���S�P�>Z��˧�46N�?i�IR�}�R�`��Fr�6�to",�8\����?��纐=3�k���y}��*$䵗����#�Ǔ'�5�d����8���W��)ݥ���ѼSJ��aGx��Ir,ED;�����I���C��7�X�����W��.Bˮ����b����T/d��rp���t�;U|\_/���� ;A��cc`��GeR.A�ov��d�y�)vH�Fiz׽DK�D����L���i�pi:�q�ϟ?�J���yOV������2�E��T(CP�7�Z���Ozj�������Q�
 ������=M��Sݝ2Yy��]���j,�Ǐ��>�>�w�{��L�^N�nk�F.9B��= ؘ���↘�|ܶ�k��F��u'�k�V�[��f�'�$m\(��`�m<�%t���B�{03�_U&�8.��h�A�� Y�ˀv81�z�<�(���}cƺ�QZ����֤���T�yӳ��J�Td���gxcdw"VXNN��ǟ��b/�?��R{��O�ёǽQ�‍���Q� 	T�T���;(r�c���� ?Y0[.T��%��1�t��e��Hz:��QC�_��ͳ���0�wZZk�I:5���o�T�XYX`�����U���߫�t��%�GMe�Wl9^�|�5���!�����Ru7m2�)�&ks���+�Q�<t�����6�(7d�A��1�����+t�ur��m
��W;�����|�{���� ����_f�wn�}�!��/(@ڨd
�k$��()aifw{X���V� �av��xh�%m���P<����`�B�l���<���>���kk��z[�M�x��{n/8N��\\j�[�p����rb`����R7o���'|]�.X�m�nШ.]�TdMN��Vo���u�O�g>��/����4e/����q�e�_�n�|�o��R����'�Z�K�͚�򌠂�	�p4�����_��,�K ��$H���e�V��k���!����	)LԾ�U?i�hC��MU�y�
4�bׅ qppTl�L��S��.��#���Q
�_Y_+t54x�+����������5h�PHa�9�9i�󺻀��`Q6��ဖ@",���_ c7j!uss�zt��h��@"bϚ��Ӏ�N�����v�$|����O��vs2����̚�fC6C�:��\x<���s���|p�ͤ��F\LDfu2���"��P�]zHW2X�(��_I6Aw���p��ap�
�v4�|MO\'u�]H��~q6)�Ŋ!ٺ�9N}�B���O���"_)�A�n�B�.�肵}715�ݽ�h&��F��,�<���� ��9Jlr��|h�I �;n��Ov��?5�d��'� ~�DAE��M�$� '������E����� q���"H�T��c����͗o^�*��Pq��[�Io7���Up6'%���')l8'�fWSCEC6񾰰��P\�4������x���yCw𥚎}(�3��1�.�����m��I��cq�	�g��D�H�o�om�3��e��#�T���M��*��B�N4��ݯb%.��[�^WU�AH� 6C���`gi��	�s�ϝm�U�c[�A�6! L;����1��+~tC�:�J�����*Pd�? �Ԅ�>ָ���1{˯��0� +�O������B+�Tw�����\YN�髁�g����C������,������:aH��!/,.j��y���b�����I/zȌ�'�۱7M�b����%5Eǹ�ǹy��Ff�[$��>'��DҒM�o��(>��o�/��Z+I�\>K�/�O)��+ȱ�$��W{ �e�\nm8ɿ���E���T(���w��,^ ����h�I�Hgam-!Q��3���e���-,?�~g�{ f`� �Ė���o�?��Z��P��~�Ȑ��aS���bHB#F�N�^�Ȱ�L�E�.����M3LA���`��L {t�"�[B��{�(�n� 
��a�"����]H/�p5\��'�mE�L�uS0��h��`�u�BT��Ŵiٲ�r���Th�1�d�c#�pk:#�&H � E\��\�(�N>0f��?� .o�كOlVÝ;}�5"_m�q���B�ؙ�~��T�a����K�z1S�������Y���y��-�l�֋>���?8��gB�n�D+�cɀ��6iИB<J���[�w*�&dX(���z�g��U��'-��>�f2�.���"������.|����0�0k`�N�	h���ð�������MOO��٢aF�6
���ű��6E��1z|�����?M�络ɀ��O[\f�`�:ۆh9�x�Q�`�g��2�!��}N�4�F:
�:��z_ZzW�콼�yh�ye������n�Y��} +x���T �.ŶhhkG�Đt�^� ���t0->�\{�D�x%��6�@-T>���ewP�����'c�?��//I2���pt*�:���3�K2��(�{pၐY��QI$�X�{��^Ө�}^�t����211�+Ӯ�7�ɝJ>x�����J�G~����C���{A$N�жz^���`gT�cW�����χ�'��(_� �*2r���,��� d�M~��_�<W�Zuf�!kG��zR��uz��5�x�&�O�p����u��ʊ�>)2T���+~��7�� �;�1�z�2Y,(��3��4-Ez�2;!��Ͼކ`�|�Y���C�v���og9��y�s�,uaf ��;�͘c�q�\�Ď��ǂ�$��H�M�Ae�Zq�s��z�꾧���p�U��SV:$@U�쪾��[��Z��ӧ�OC��L_7r������d�����|-��?��{ÿ[�KC||p9����Z#�o�\��	w��:�XV�<�O �f:�j���&�<��L�,�
n����6��K�
+�-Bm�8lϜy���nֈ�.I@NC��;F��W_�a�E_�����dN�Wqr�8��Zq��wvb���֓L�A�mVz��C�H�������#~P�ٽS��;�cY�%��v����T*��$�מ���t��O�Io9�0��{[L�����)Pʐ�q}��������T.���M�i�k������	,����48
�$7��F��&}?��g�`�$Ӈ�N(�3���F?{#	m�&�G�Q�/��w�o�~���
��Q��Er;���1�M�$iiY*K`cm-el�d�Z`�dfG&���uG�2d�,���&�P�ĸ�_��N�Y��A\��`�̘�l����x�z5z.WDDĴI����Q�h(!iPjm�_����@l,HQx��6ĩ�g) ��W@I+)nr��Nj=?=&O�����嗕͘��H��13��0N�B��Us�K0pE�����oya *� ��#�E��N�g������M��e��{&0�H 2���i�N���S�U�fl��^��;aA����ѽZ�DzY�H&��[��h�Íd
�'� .
�R���ihh�P���p|ײ��vj���=Tl �����^�_�͖
�l��wA�>PQg�2l)�rɟv�u8���O+�އ5s�h�:�D\�2,�VE�ۭ���0�V�PN�ل����X��8�&g���iK������uu%7C����XE;Jr��?{�f}յr]=&�z�
�� /0�����W}�L6��� ��q�6~	�А�[|�P�����Jtm���Y��Z|����`�:��.WU�y����V���0�Z%��Ԩ#�\�C#7�������� �v�rc�`�{>56�ӽ��O҆5_�������塚~�|)�����vL?�^��(ϟ��>�Z�I��ٳ�IU|��I,9��%B ֊ҍ�j�ćJ���o�oNM��p"4޾5ӣ9Y�Vaē��gχ9���b��OL��k[�]�uL���n-!L��'S���HK��5�=��=�# q:yT�h4rA������r'��΍��U��l���"�8���!�����9��qN�8�kh?�+���g��K�nԔ,�O���HO_m�~D�����͛-�N��_PP�?^����d3v��y{(���}q̒���ɠ�����c&��z�4$<4�����|L�󔶷��1����2c�[��E����������t��?�қ�n޴,6�G�V-�	�P�0��q�;kI�;����~�f�`���$�Q��\��߹d^��k��K�Q�pU�kkk�\:� ��A��&	1��x�`���&���O����W�Ũq�mMf�֟b�1�(��k��z0�B|���#p�6.�_�=:�i񺠔��G�������A�6⹸����X��6>K��Z�U�K��0�֊�Qgz�&6J�lU���S�L�v\,����dIX�}��=�`������t.�YǙ�� �m
��v�F^[��<�X��Ko�]8�P�Ї�1�1T2M��o|O��1�o�=�BP'j]+��y�`7�T(��T��7qtTT`���rB��^�e�[����P:Z��ckN�_$���.7v�?�^�K��� # �*�:�㕝*����n��N)�܊���֙��I@�6/��^D�:�u��4j%g``�lz�m���!|. ���;���2PV�^�^�C
���!���>�LZOa�A�;p {����ūsJ��� �#>\�Z���PEN���u�<��×�^=�5�g�	*_�M{��^�P��C �0�?�>�Gkyɹ�fM/.Ƭ���'B����2���8����c��3�wGxd��4c>���N)��߼��� ".&����,̩��F��J��<L�"s|��f���l��N���r�_�{{{{��:5[A6p23ix�e���eq�p��w���+�,�Ep'\������A{Δ���:tt�Q�H�� �:~%�Ҏ�!��@�Ѻ��	�?'��_b��IT�N��~J�l��y.����r�B� V�2����" >�ޗ W�t*+�W����z��xC3���R��k�ߚ��A��zl(�R�l��&?�:�!�=Ի�J�'|@ť���nە�'(o)���O�K'"^[�o+'��X�65�}-~�(��@��u��/�텽��L)�O�=��8Oy�ǉ�O���I5ޖ�osLĞ���ݔ���]	@�x!N��b������Yv���"=%��f��E��jI;O@��K#���8�e�;x�p�K��ï
���+q:Yt8�@P�Г!\C��k�R� ���K����p������UW�����ٙ���f�I�uG�11(�(l�0�zyy9C����]�ϟ?zN�@S?�����>ۊ~>	����RB-O���29�����xo���akz�������F��Pk�_ �4��3�f	�qǬG�J����h��1HI�0E�4�X�L.�f�p2�G��&%'�JQ���y���=�U�jط����x]Cø���əX[��	�Ҙ��qt+!A�y��)�Dɪ�1���s�;�_~��N|EJ|^
P����j3i������Y|pLp)�g@|��~
�-�<��>*���)96�Pu8Y8�u�l��A4�׺Uh�Ʋ�g
��D�r���Դ hǭ.UqO�N�?L�;��RC������)��j�Ԑ�Ⱦ���>
"9���d�<�h<�ܱ�p7�*B�jI&�Io@�;�%�:\��$)"a�'&~�fec�6��I��y >��[���p��������H�����?�������F+�;K�	1��M?����c�: �*��?s�s $))M�0_oG�y���ǏZlcTʪ�5�(�5�Z��!�~�#eg`>bW�>Cx���/ڧ��8+˽=��g>T@tgt�h�~+(@�uT����gn�t
	�r~~b��>�u�޽�k���g!���(��^>�Y(��8��t&�<��2�D3B��jI"��W�o�u�����m�f�"��
|<::Zv϶x���j_]�I7M1%�#���ę���DY���ޢ�Y�=R�������������}�+�V=�{%I��=��������J��ᣝ��8���	���t�_�hղh�BX�fpW�[���Gm�I�3ƒ�mr��Y�U��XW����W�� ����N)׬o}��f���X�~����H�K����B�h��0$��R�W��Ot�G[�b��g���؏t�9غ��PX#2���ٗ��\�&�k�J???W�Q�4�����I%�}z���ǒ����v!�Td&���(�F!Z����..|����֑���O���X(I�/i������+�SJ��r�]�?U�wr"a'6�WN��&�H���~��	���\{"���?�����_�:�Y���Җ.����h��a{�ژ��� �y�����옓���mo�䫫)� B��խ�T�όe�>�c�a��vd������ �q��נ!��엫���8�p9DҶ�=f]�6�['8��3D�*��^��=p�/�0�to�㋥|�b%��H���pQGe)P�~���= U�dC ���<񰱱!�[���0ѵ��1��7������-��;2֠�a�ЋɆ�� >��~�A��[���T��jHv��(�c�)�&��KA)�����k$~(�����>lm��6�[����p2Ӂ?������HM.�߿���Cp>�R?�� 7�[��P˚�#��>�]�X���	Ϸ�#��/x����.ӊz�����B�߽:WA�q�aPǮ�q�bwsy<ୂvZq0F~f���'5�����c�B�����I4��?�3'JG̺�[Q�A��a	��)伥n6}ju�V��"��$�kě8S�v�0�vkk�d��?V<���M [NB�Ԋ����͉��;6�v����ǍC����71"�So�ѻw�6^��:��3�I���-�@��K��H����txq�N�sՓ3�p?������r��\/o�
`@icgg7��O���V0F���@� �P4[^_?�t�77���� �4)�����Ծ�ǽ@G{���SS��'�v^��G���.t����B�[�^�@_��|��Y����`���/F�O�Cx3�欢UG�ĥe͞��̴��WaLƢapXX�X$��Q�XNت����)&��eE�é����9���M=T���΍��Iy��`��	A���k��f�i�op�&�Jo��	��F�(qܞ�l��D�8���j�C]:Y)���f8_��L�1;+�/�0vw#�d�����Q�B��ߒ�j�t�$�����tZ�n����{{�/���ǀv"""؍i���7��͑Hp�?.��PJB�j9.`�h;��0%�7* 1GJ�J��Xsb��NƉ�����_wL���1��c�|'_&BU_���,�X֤�FMk�/"/��kt�teD񊚷\��_r�\3� )_��Y�[P0\��5�����rOc�M@�2�� �+���ߖ7G����-�_b����m6�͇��,u�(�ǂV/�����UK��
xA�ݾ3�S��7/	�̬��3zB�,��7���17� ��%��h�iu����ܼ.�:�q�{mB�~/1�@
T���HZ;�E��lt*�<����ĹOJeҴ�\�
�h�!+����=E�����Y���Y��q�sų�&����}�g	ކ܎"vz���3����jfD���5�"ʺ/B����%����d�n:���NL���:
���7����+-���-*hNB�Cpm���
^ 2F~�~����Z�������M$���q�@_'K�H�(��0b�'�Ѿ��|�΢f~rf���z��K��4[�I{���ݓ�co���\�i��!�7mkT[0��@.Ƣ�3eY�N���h)���2�n�,�ǝV�w]�b���0�	�4��`�	Q�����efv6���@l�x��C�U�Eյۡ;�Q���NAZ:E@�a@@JJ:�i)�n�����S������w/?��̙a~{=ϳ����g�U4/�t��e����6X����Ѫ"_�E�KJ�Iu�t�oP�i,�K�Ͳ��#�بʨю��^���t35d��|%~F��[��Ǖ�e���Ҏ?�B\hx3�MdoO<�!ea��)otv�u��ʧ�#;M�l;�,�K����˦�r9%���p+E6� ��1	\9+�Ayt55���o߾���_;�����T�S�9,�4��]fB.���@��Lkn���Xy ��}$�gy"�L�4�pO�of����˹�y!���Bo1��'�����JJ|��!T����#����"�o�*U��l���$�e�G���Y���,�qRĐhB���W��9{�9�@����Ê���.YG�╈],5��;;;��bәb)���?~�E��>4���,����2�ߧ��>�ub��B� ��
cXD�%�E�9�%�3��3L~<c,�	�ktʖ�(��拯��&Ya�A�vO����BV.��H7j+��[�Aʼ��O�[�,��U��ͳXmW����sk���k<����'ξ:��3O`@�`�B֛	��M<����̵H.$�"�^�*���B����rXTʹ�V-���`2&<{�/���l)#�)C��k*�_{َ�g��P �mh�N�&t�S�>��mP��@�����D`hd�82&cd4�s�}���Wx�7�䐐ɦ���i�O<�BN�����
����}i�3]��O��w�NP�W��K[�E` �'�m�M�ˍ�0�}Q{�$(	����S��)O ��Y͸A����$6˧�t�z������@�yv:�$�k�f�&�&I�j���:/����������dz7{J�����������~�i���Eq�E�\�pQ�6�ĺ ���p}��ל���û����V-d��IBA�h��Y��wc�}��؃�V����$OV5�-�2�%m$hW��C�zTQ��1�/�Pl㮛A��G����m�o�	^��^�x]���&�;"�P����X5�8�wO�!� �;CCC��rk�k��TL��r��9���].�-:�j����Z/7��R$)�@���g��U��̳|n�g1��פ����s�,�|r"��wx���*�O-�*��:�c�=[gOΐ�xUPYISm�����>���/tG��U��y�,~�0W�G|�/��*�2D&7>L�c:��lw��iQԲ&+`�\K��]y�ryE��7鯬�YW��WEAc(!ad�(�y�)f��+��`��e�Y�E��P���w���Qըh��E?Ǥ�šwR�8�>��j�E��C����X���Ag�&9�Uߟ+jC�I��z���mQ�V�I}5b��9��v{�����m�����(�go�6n���G�ńk���6���r�Ƴ|��UO��bs�Ȝw�?�/��G)4��
�b,K���o�4q	������J;5Ʀ*�����@��nft$C$i�4|w���29>Nf������5G�a����v����˩�����S5�l>��a%Vr�7��W��dr��[l6��փ5k��J$Ux˚V����߻��H���k�mʂ:8�1x��V@�N��%9�?4C~7K>��f�GV��E�PG���A5$��U~HD�����rE�FUh̛mf!Qy!"�x��IϘ���Cj�Kxr�io�!IY�ɐ��F��D�G����7��<��|m̊3�&�Ѵ1j�b|&*2фpey9���5��K^��E���h�(d��9���р���º�T����c�<�o��$�(Vy�ǘ�++y�nM�^�k��pKR*�[>Y�����Qؙ��>Bx��3�M^�J�=�+��݌�둌�z�����E��R!q��Ҍ[H��i�y����z/� �B)Nc^ � 2@�a��1��=A�(��٬,n�}<�{�����j²d&&&նUm���$����W�3�:J��c!�V��,�6�EI6㻟��X�|�J�a��::� E������6 �:2j���QF�Z����~O�?�5�3�p�mC���]�T�ݔ��Ί���gqJ�����a�އ���_��������C����k��n���P���_�KE�Ҷ6	�G�Fq��3��U&�]h���X7�5�_�ݲ�)���[9��� I�L��d��
p^Y�����!eb�I���"_Q�����,�΁#��w� Lyk�n[Lݬ[y�7F�|�|3�[��P@qL��/������&=[��_?��l`��I2E��'ě*�e�@g��;��m��m���2�K���J����!Q �����kFYN2_n�(Od}��5V�����%�Tп*��^dUc��ȭ���?LR��;�'t�����>U����NV1s�b^�9��v���������Gd0�����j��"ҙ��#z�ȇc]u��s꧗X(1�$$Zlv^�zT��:Hf����~�n�q�Ph����?Un��E�IT��m~�SG�����R����W�n��wC�K��R�q����q֓�� ���Ӕ�k*�b����������A�����qׯ������U���V���v���-)���C�v��m��>��tG2��"F�{��Rbg��:��gL�[���r ](����[�uo������Sb��/�8��r2mlKqÀ�1YT/��^�pzydTT���Wiuӳrx��P��2���>�x�nM1w�b[^Q1z�G���U�~$!'�����9�ALY_{������[�*�fKT��q���M�o�&��n��bw��{�nڲPI�|�n1��3�[�u�.���o�_ܴ2?f�d~*���[t� �D��>M/1@���B	���A>��`���*���}�A!�1��x�|5dgs�Dp@�,��������,��;�}a*'{gg3F(n���9Q�z�B�Q;|��艐�Z�e��-Y��*�T�A+P����m��Q������5����߿⦶ō.c�qc� Ѫ����}#�<*�>[���0lu�4�����٪_��./�����)Oi�ٯ���6[ﱗ�i���hDm�	m*��K�%�,�d��3�,�=��o��m�}�L�D �T�;�*�1�oa��U�����^�hZ)�� ��9�@�����-s��o��2_#q��y�1�����$�4y����{�b��0��Z�7n�x��4���<kr�v���xG�b7���"�B�/�L@>+���#���GN<�D�*Z�)�W�h��?j�8�c�233)�N��F�$�	xZ�AM3}PaH����>�b�����&I��s^);�����.輄�=�U0��y�,�ɪ� o�立��a)�Ksˌג#+uDŗC����� 6�?DZ�m�29%%��^�}�7��^�^e���t�۪YNQʒzz,����U�d�vYC.��RA6����b���  l]�	`��APdh��]�K k'����������i�y����@�sTw��%s���Y�*Ǯ�����I���f����]'@��j���߱u�M���*<��X� �!á�J���Z��HL��Ynt�(�#v
������H�f�LNM]��;�^\��{J�X����w
���}���{���cғ>wt ��Ϗ���=-����1,Z������������7�j_Mܐ?��/<��SZ��,����I��=
����7Ui�@�X��`�U9'_ �{�=yYyH�CU�8$A��76��N��4�9A}�Q�"�q���s 9̙�;�%�OwP��xz���o��]�N���Wa���A<�q����-")s�����v��g��KxO�@�V��f�B�.���Q�s#��:9���.����\�S�Aƨr����g%�������4ȵ%"����7���"3�?j����-�M���wY���y�?�IA�ʕ���苾ڇ��wkg��{+�{��I���~xs�^���~�)�e�;U;;8��:;:�V[�>z��t�<�����+������,�Xm�)GTא�����ӌ׋�qQ|��`fy!�<KA�{���@ӱ�4��"`�7\T�.$�z�T��o��|��SQ1�2�f�N����iR�_�ψ�-��͋>���H�����~0vU�QHD����-,�h� �&�<�+r�V��c.���Px�O)?}�i��*d �qk��-�p�a�V	("s�{J��'�x���kB<�:��@�5t���5��f�����<�?M��\�D!�v|��� ��a�sވ�\�/�ݑ���S4"q�P	)�j�S�N4r��0�����>bu1����~	���GA?� �sD�W}��<~���TA��z��x~�aE������� ��W���mm�$*���/��S��ކ��
 �錏��`4<�&pf�[[;�����ގ9'~�z����pm0n���W�LQ������"�61�W)/k��Բ��:��9`1,��t�D{�U*MRP�C!�k2ﲛ+��N̩q~rV���q��%�(Ѵ�d��=wtw�jrA�c�Ru��) *u�pwFS_�9avt�>��dn�?k%�������]���y�XM_m��Տ&����ϳ�WL�e:3�Y��S�ٖ���A�,t���[D��s���Kq�"���Sn�5rG��9w�ƒ��-%����K(9.Q#�O�.��D罭W��6ӕ؃L���hUV��o�n�X��$3B[�]*��=�Bܪ+mYZ�_�6�b<c�ŁRAQѪ���9��M�"����@w�v�Y&p24Z��M����!���;�bG�Ż
N��W��o��e�b�������3�MM��
3O�G�%i�K������.����z}f�r�U��0Ta_ ��U��ؓf-�Gl�c�'����l\��68���?���%v3V�l(%a�ڂyc{\NE�Ԓ��^�lp�	�Yw��f�Y���ً�l�e ����Wr60�F�i��I��M������Io�K��v`������M�`v���̇���>����_��f$;�p�T�P�1�\���jlg0q�6k��X���&�9���$X��G���Q�KEl~+0�]6�)b���j 7����hKJK���?j��z��RY�*��az�8cpgzH��޶�����Ȅ�آ���Q��*̎���I����AL	{���+>�z�}���r|���ޯ�	#7a����WĿi� ��DuD�!`�j}�B�RQ�?.U�d�@����LlΓi>��⚡�Ƃ�������y7��'�*�F� ���o��%q��? Y�o�����&5N�^]YY�z���+�:$#���,�ϸ��h����د�zߩ�M�2
�v?��+��i˼���F=	
�_}2�g�y�d�������i{�g���\���D�����;�Vػ��k�%e���on4��\)���m����Z������h��6��P)k=M� ��������Dc~QQl��"tK�̯�x���rE��>NW&oФ��2�A�Z&s"�VG�w0� ��� 8pR�AwP՞(&�ӿ��_ۤ@ÁmY��N��2::����s����5L���\u����2��QS?9��˽·S���v{?��[nv��Xgy��A��=��`d,��}$5t���jc���tt3�c���Te(p��)O+He�X�B̗�]���d0�o���a���B`1p���[&��
��V���a��R��k/UU�Z��ᤌ;�X{��e8{�1��{���DE~4�VMM�$������TyM9j�=n��ݥ�ߢX�}��\��_R�sh�ْ= 3�
���9f	��;(��Zm+q�a�m7r��ˮEp�X^\�7y�Do��5��Kuˇ���^B66�Q'��xo�}�#�͟^Cj�!��=����J?�E�o���]ۀ�#���F�I�&a��\$ع�i%��WC3������RI�5]H�e�`Q����z����kb�K=/}}y6xw�h���WSl½�,�����I��lllA���E�(>����yZ�Q~jj�1�w���,H5��f=tuj�{�v7k��h�&TH�l��'����:<×��?���y�ȯ��;�*��Y-)!
�������ТD�a�n���(0$$)�W[�T�>���=��̹�8/M=�e��8�uK�P"N{ �74~�_E2�^��l�>��!4j��|ĲR��B��z[�&��2ss�*a�K������ � ��Ms>��qok˶�E%���U�#����w�]�%��OγWVo��Rw��$�?s;�U��!���sk�����yVE*�I�����..��?
u��0U��o����2��,�����& ���uR��&ft��ԭ�����:D�	�6"d_f!Ý���ܼ�}ie2<�QgV)=���3�)$m�����G�:���&��R��C�[o|�ī�y#�SPrbp�C�����	O�R�CܺKtJ���3�3��5�����U[�4�Gؖ��(�$.h#.Ƌ̖&v�5���s:�$L�≊�N�?{�D��͹/��qy��E�����ތH'��6Ӕ�%����8�	-T����$|�Dܺ��,�����,��" e����SeU���Ln�uә���O��imjV�Ԟ8���v&{�s��x����%��;�J����L�3�����P�x�~��/C���B�&�};����C�N��US�#~���@���S����ߪ�n>�suR�gV��W��a�9E����i�i� �ҪO_噿Y�x]
�7��g �x�u]a���}�z���egwMZZ׎�"��ԏjT��s�s\�>�++t�FFV��c2��;�Z�^:����8c*�,p��S�6h��PZф�V8+q��u�j��D�i���R1��� ;v�%�c�j�����Ԧ�ȯ�T�+��.��!��[�e��ᮽ�W���An^�:����<�-fv��\�	ڗ?1�{zx8 �<�tF�w�U*V�W���h������w��X�"$��s��vٝ+n���g��jy�ʕD��FY�ZQ՞�!kt���w(6azhh�e%��
NZ�=��|AQcͣs������hF0wɐ�#	�A
�q�"�W��@Lp��*%�J��0))il֗�:��T�GjOOS��YI���y��#t��H��I�49��Oߡ{���5X�8C)��f���GR�L�w0q�E�����h���\4q�������`jj$-�/r�rT&S���u��5��A���a��x��4q�ɠ���hn��G��;�|	���7����aJ�s�����'�ݷ�@�6E�S1s�Xbm��/Y����7::��$��������,j0֜�yxP^^��n"�v@�(��wݣ$1$F�V�u�_痮6Sl��_b-n�����!/^J����0Qd�PY��_��]|�]���b
�W5�A��'I�wy��R��J�s��O7U�pcJ��q>�ӿn�B�f�I6���Q�5���\K���%�Q��Q�]��|��F�F�� ��yQ5�Mc �o��gb�����'��qk�ed�sENUY pxZ�a$���G>Q`��}ծZ�"�Ч� Xߥ��P5���q�'�p\@�k���)N���w��Q:=tx��ʶ�w�W._�Xyx��
�C�^�A�HUg?�s�$��"�Ξi�nb��KQ�]�d��"r�-��]�(9!��?'���4%q~oNĚ? ��j+��^\6Ɓ $�"S�5,b�o�r	d��i�x�H&�0��t���0�b��2Gȅ�C��%�7H��`F��6��|���}�ԟHN���ST����L9G`��G�p3X)����j�h�f��n_-((�-���0�?}�e�"�����_��x���W��ͦ蝍��n���lBi�{��qZ�݊gk���i���%��������.���33~z��6y�b�EH����=i(���c~	���t� ��i�%	�Bf��b�[�|�:���݇��t��&7���XT��[��\���(��B�ce]���J+ ƪ�N����S��2�^4�q/�޳���ظ�z���Y�a;Z��'oY�f���퉉��_���~��N��Dǖ�+��g�Ǚ���P��<R{�&v,����C�%KR�l��K�Y�a��tВei�T�����[�����wR&����!J�l+����
X��Q�*�����s�S�c����#`yy�Oi`L���R�
M����V�h�H��Ev�̢�X��!�����m��s��VkuF��	�=c|�-bu4�>�*4y�&QM��DH�>+R[����^KL"^@�Ҏ�_&���U:��G=���]�
�h"����}�O��,��q���~O��Y?4#�9�2L�f?�E���S}�T�	�é~���-���p�1�]����7�"OY�2�᮳ �dZ-
��U�� )4r�ve��!�Ѱ�?	&*/t���8�e�Z<���<�A굱�fNժ�����c��,�|���N�Y>*�-�G&Ӫ�U�y�E��W$g��0& nq�E<��e�ϐط׃�D^�K�T��k=������Y���@�r�A*�^��� �����EJ��;�Å�͊���e��}�_:!�w%�]�gr��.�l
����~T 
�����ی�H��V������'D�ǒ8�V2��!�Y��F0��bm�9��1d���Ox��3-���t�x�U�W](��>H{��*��,}�"C*S�;���.�{y�aܜ����k/H*�|���r��@�KW�9IZ�HV>�"Ǿ������TA���c�#{ۚ�A)�Y��߾Yg�B���uwU;d��M�c��[�h�*�t;�;�M�`�p���S� Y_�!pJ�@��������=*�z���;�� ����q?��nH6U�Gxnn�2�ά���
K�.,��[�T�h�z\�P̻�7��E��k
����s�H��ي1���Z�&%6~��G����x;���[��r�fw��c�ج!!tu91f��JO9��H_?�Z�-Y��|/��[��F,��1]��F.��	���P���!@���I�����n�����ÿ�b����>_���8Yɱ���u�e�]t�l�����f��9Ӳ�"�����P���p�cr����|��Qq�5r�l��{�ƞ���!��+�`�b��6���a	<ß���mf0��r�<�����Ra�t�H�8N����aF(s� }J%�Ye�����60(ׁf������cУJ\��PH��̋$��T妚����k�A�t|.��Q�h���ꕀ��pl��FO���U�f���3�4�����	0�Ҥ �>�B��$9MOG��ϟ��ҧL	Or�9��le���Y�#����3I>9�՚8�	;�����R��3G�u��Z����s��m��aɑ�	F���T���Z o�W���n��}V� ߹o#�J\�j"mk��6�%G���bG�w��J�EFXb��͛v�[@�cng߰ͲE�k	��[v�>��g�}'>�����n�O;vv�|5Q���a�$��Ɠ���RQc4�j�蒱8V��ҀQ�bj�$����4F��5ɹ���Ꞻ�)���/??#���ӧ8N�m1������~.m+��{'�O��8�a�u���M1�N����BSR�=�}�Z~G��-�nӒǓՌ3�;���tP����:��8i��#��uu�,�5�f�3r�Y �Eb7;������B�!�}��N谏Mx6�p�(-$���z�If�G��|�44D�I�@�82�px��m1$�H�Ơ׊�U��3tJ���A�Q�xbW����S6U��8ΎvZ'���o2�������L썋pth(ڬ�@7rd�Px��X����y�J�{�~���3S�:��Z���F[��O59<�;�5���?g[t��o��$S[�r��3#�9��t�>>>��W��zb��J^Sβ0�f�I�$�6�i�:���o�~�Jb��A��~!mg_ ��a�^%M�QuM��F�l	��9��R�.^�V��q+�^��:1�Y����`�z3&.�Mf��Ɨ�����^^���h��R�kܗ�gR,$������P�iƊZuՂ���`��!�
�.���z� �� ���{k�s���^���iD�k�\n�#�������h����{��
�> h���!�<��U4s����2����A7���9�}>_���
x����%����eޓ�:�v/��^D�a.�VUU���O}�0����_�Z��l��U��󋋘��?V��Fv��T��{?N�Z�`�L�<��FO�46O��·�PaT��io�=>>��T$ ������h��\?/Y;�k{q��F>��1��9=��P�eӟ�\B�cY��l�T�h=�]�L�6��ԇ����/W:�8��҇|z�\`���j����yVm��mN�G��Y�ܳ��# (=gEzK��z��z����M��9zV\�>�D�
3 ���N�%���%ϦS�Ģ�'���B�ES�8�ܬz���uu:0���G��������>��I,�/���ާ�'Q��U �jaa�J?�Eݞe2�O0ߡ	�ڗY��Ɵ�,��c�(��#%�xA���+2ss���`�&�c��P�h�(^��6$������������^)>���_���oJ�P��U�a��ˡu,��VԪ�Ǫ+l��9�V��BM��--�0ahh�r�&�o�g;ɋ;�H�~b��ΐH�~*�7/�]zf���gIp
e}����@�L�|���.�)\|�#W�o1>I ��,T��]\Dұ���0����C���v��/y���vUǴ�l�j�~��L��"ɒg�7�0���ec�;�v�+�2��F+F��G�o�m4�]� ���7�����|8ݠll�hى\%&�%�f{�+E��7��Q�N�����dݷ�z�R���2�-�A�
�T�S�(�ϟ��7u�EmY$��]>_Q�t�%Q_q%+/�⮛lu���ڀ0��%�mpe8�C�����k�E�3U޴�|������m����D��A�Pi����Q�'�������ۤj�\�����<�����
"��$̄n�(�fZ�q��2�6�S��L·�.��5`���BjZ���k �jl���o'|4`$y�� NOV��7%1��!�O��~c3℞a.� �
��)�Sⴽ���M��ܷVa�����;kt̘�p����7~����)�/�k���QK��S|%nh��dEr�����ڝ�@���cI2슸���`�FW���k�ܙ�W�>�5�w�x�9�����!�h�s�=�A��~�1w���&��)2r���~��E�=	�(y����uɐ�%*�ʊ|�XI��,�ǧ��=D˯<|�tA�������;ۼPלge�Y�ֶ��P�_�d�}��G����Rµ����[V(�&{r��U5Eؓ��o�8�.f�=,ə�}f�����	�^������i�U�+���A}"_��ns�
K鷬���N9�dQ���層�����wF�����a����U��15�<�mX��l_#t�6�{ϰg�Q!T�e�N[婶K;b�'##����٩�CT0������KnV�{B޼�L�ѐ:��r �ֿ������ݰ��H%�@���8�d�fZ�
P��+Ziܗt�� ��1Y��LG��� ��whoԕs�-}b��%��TN"W�j?nH�	�]��i�SE��~�H��ϥ�����fO�!9��q��x�0�ŗ�+�������>�U������H�ܡ5����cP
��q���lw������2ӆ�B1t�򦥥�m�������S�H)B�p����/0�}�W��	K�&̆;p����& ��a�����}��x-�����
�6��3�^
B��ė���ո0���� ���F�?���@����_iQ�M9]���T＜Bݭ�V(=�˖���4|j�-t���VS��p8��w�a߃��g�M #z^L=���aq,��l+���dw���;m;T����,������;.����a��ϑt{�fA5]_,��n�a�V=�*=�C� ��k�Z	H��Fԓ�(�~��LB߳��\N���
ߪ�~�]�|~�z������W�=Πߑ��e�]�M�~���S;[�����r����$P~�@��f#�*�s:�r0p���Dţ�3�����ʄ*�^��'[�D��N�=�WX�1_�,�y��v42�b���Ț'�Jv��7��8��/���jEV��qO����xL2.444��u������i�M�������Ɏ$��iXt�_�b�H��D..�k#�"p��&�@�F���ݼ���pM��K�����@���c�O��ԧ;�I&8����d
051��P��(�^�Lg˧_�d���1��2�yR�D2B�^'O]�ŗ�/E���GA\{�]g�>~�Yq�Y���f�|�u%���K?�tO��Ǝ������M��~������]Yht����j�v�o�ib3��!I9Py���5��W3��� J�,�:�S�E�U�,�n\K1�ӭ���=���X� m�:}�Iv�W)�]���#�@�E����ox�&����F33��&''u��K�I�+��t\�e47"Ky�˓+Y���j^EB�S���5ٓ���9@lW](��<������%j����Z���q߳���u��Ũ�ҰS�3ޏA�-����;�!��5�k�q%ǟ%���O&z.M"�.}���'�
$Z �A
��1z.��{�Ά� ��*�,Z�@� ��@G�ߧ��aYD�73�͓�)�����˝�.Yww~��nZۨ'_�[�
�j�62YL��CV�%��
��FG���źo����1�--}
�e���!O����r��E��eG���}4�z��b��zgډ_�ɑ�'��T�2H��{^|||��ٓ#_F�R��]p���/�X���#�x�x@�~卮�&3!�Ͷf!)}O{b�Wm7(✇��SR2;�<P���J|Еb�Tr�/� C�QOՇb�N�w�!�<�?� �h��^�^�ġ�sMmcK����(yh�E~��X��*3����b+̉��	�k?��P����N��P��'�'I={F���0��8��!�%F��3�跀�'�w��tٓى,D[\��[�~�ߐ��O)��*�!�h�b9>��sK��V�������y��`�y���k���8������Q�<%�)Wo[N��k�z�����=�[,�В�,,���'��,�\�m>�kO��]WHP0L�������Ϟ;��R�|����&֜?��BE[�,|��PVT�z-fx������p4d��IJ-~�#BӼ�q�n��M��i@�U�]��9����ؐ�����k������sS��������h��m�cc?��j�#����@z��j_Dސ��I�Ƅ�K��	�%Be�\�7} �,4�"FY�X[ki�ag����Xx��-]ʻ[pr/z����94����Ԛ�s�/��L��&3_����T�5_wc�n K�p�N�n���`!7��m��|������mɝp�s�����ߕĔ� I[�89�$R��
1M��ם�gR	��`�a���9ŭ)�j���|��weɋ8�-v�3_���z3��X��NNj@Bۦ���*��`��k�����
��:!E��?�@��\y��v��-�	X�-�/^O�ۿS+��=w����:*4���^&�h�St*'���ziAO��2Se����B�U!'�^g�W<+�%�.�]1��<̃}Y��#/�m0�@�U
�ȭ��q�C�2�w-0#į�ڟw���H�,�k��*�nn�n��U�n�Yf V�'P���'���AA�ԩ܂4���/p
{��\۳�����m�+ZaGd����b����F�-��"����j�'L!R�/���m��g���;ԟ��mj�O^���\b)���ﯢossCx	'O@�d%�jpߊ�,�7��5)�_{�ް�}BGw���B�(�>����{����{@E������0p���]p0v��m��s�
=���e����H ���<&�g�d0�|��%��|d���e1���ON2+���o���l��g�8ȣvŚu�17�tll|Vjq���TUUA�X��#����D}Y�`�t+K�g2�s߿�t=�2��`�������)����:b�	LT�M7D-�}��@�������AR�u��KNn��4��?�%�+��/�y"�P�Bg\�v(�7C,zЙn�dD?{�]W�R��,�PU@H�N(�cE榮 Ӊǧ��`��9-һ���2Ymk^q1Ve�Y��q�D6����rA%ٌ�Q�Pש�����,��B��5��9���^���L.��G��B���d&_����C��J�xye���S�=?����9���|N(�ǘ4��J_͋���X��j��}����w �N�����d�JFFֆ�\k�������!S�I݈���C8�76��ԣYP��`�K���:���q��#V�w��k??c���)O�LZ�ﯩ���ۗ�j�����*\�����"�e�:���a��M��|a��a��t�����2�J�v�>������Q�錰�$^�'�=@L�UV �6�Q|J
٤�0U����bS����^k��ͷ&>��P�������aIN�L934�o>�®/�:3�ɀ���J��y���+�n�hI���Y�2X�����\=��RoZ�i��"=vʫ>���g�GD3��o=:��T�|ܳ_F�q��ez5��Y�@�O�G�����B=�[���X��1��q���]�,#҅"�р�ג��6�F*���ŭYߦ���	
�@$�Q��lؓ�#�ϟ�||�X�?~KG��,\`�j^�2����>��e�c���f�P(�;�E��(�}M��h��¥o�Յ�jY�Y`*��i�<�����A��A��Xv.R�j`"�9�-`JR2n-�{�^�3L����`�\c��)�<$ ���3���n��.���5
��甙�r���%�S�4�cm:a�ԈT�iX�Ȍ/�}�f�������Ĭd$.kA ��$����o���#�n��ō0_�����3j�E{v,F�o�#���ёT��_h�>>L�6���ϊ��|v�}��<�,���{���(?�M�s}<Wv���l`��0!��v��;S\XJW�7�O�&A�>����RT+<A�
�ks0��1~1ɿO&��NV�@kU����^�a�Vl*���I@@` ���Q }y����L__��jxʾ�!��ɔ�WLտr�P�F�1�f��_1��mmlm~H>�E7�@�����$N���U�R�z����_Ljx]�����n���,�]��ʌ�J����쏙�u�Aj�*}x:"ڪu�!/��f�E@ xdh����:2��d� N��!k)����(��������}ˀ�;�w�����M���iy�c]��u_��	�ps��f���w�X���[����%�v��S��ұuT����2$�@�#0]ȹ)㣄|�&b������_���=�~G��0��+!q����{o��q�sӏ$��^�R�?J������,e�Q�T&�6+���l8��`��8l7�:W�l�ً������QM��s�@�uٺ�@}�x~umF�g}�j]P؇	n8ccbV;�v��՝�y�n_��]�Jd+�_�������KC�<,n�[߷9D��X!�B�����NK�*׀Er�y�a���ק j!q�RW�m��-O� ���ei�[�QeM"��?�U\{�����8{g������F3��@	<~<+�����?��"���ׯ�q���4d>��dRZoMܖ���t�������+_�ȿ��J���i�'v��|��<��	�E��6#`�W������D��P�e?�#�Q�f{
���w6K׏�/S/=�~��~3_�*0bM�&2k���ޞ߃�V/��"����`J�ӡX�(cN2_5&C�.�`�<<N@n*���L�=�
Č�1p�h�E�h^ݼ7Z0t*	?os�Ng��G��<��4�����I�cX�����T���3Ѽ����5@�W�"�l�Գ���ɢfϖ�xq9�ӖŰ��N�l-kO'_ ż�k�[��"U�m4��N�X��u�a������| ��(��׾�8յX�aB�G?0�$/�>�涷�&+���C���dD�T���L��c�{���@H�;]R�@��^qj�=4U:�h5�_�������g�4됅v.J������� ��o��o��#a���.��(�����b���#wgj��O�wV�⤜S��e2K[�]�`�7��a�1sZe��1g�۹&���{�)f�N|�jy����"��G^}���b3����&���C�^��lDa8k��**W�|��ު�@�`�&҉83T�k�e�,B��k=ֆFF������6F�����Ͽ��T�Ԁ���A=Y��6���o��@
��C���Gñ+·pN��8ʔ��<�_0i{w��*��㞾�!u��/�>{)���1�T��u��rrU��DU�t��wr~Θ�f����x&�{g��C�O�b�
2@?�J�0N�A�X�^��s��O�]����S��.g����*��������h��B�Y�vv�O_T��;�i������B����0R�I[�o�#C3���0�ɚ�l��n^��5�G8����8콜N���?�P��,�}�������ڸq��L�3ȻW�d�x�)�h犄���#�IDC͠�k���r��jkO� �fEt��6HU��x�M�����exl��3Д��R�@�[�a��l�-Fƌ�q��6�kHZ�s�$����l2+jXntW��n�g�da�c���	]���X��5Ԝ�NE9��s�v���6�o�(�f�x� )�O2--q��ޞӲSS����ɗd9w��7#���UK:���*��7���$����/7a�:d�Q#=u���\o�𴇦<(�щ��,OO��<�=%ȯP�;����:.ʠk�niIi�AB������{�ni	A@��K$V��������y���ta���9W̜33͹�W#֞9N[&����*E��@�8�X��Z��7%j�(+������a��ʸd`n	�̓(����nB��`|>��N��u+q{�3UR4�Õ��%�9�J�x����%!�^<�:lK�?x���(����!�� f�r��:,����o�mn��f�g���D��_�A#bQD��N7���i�y��������x�:�����b%i dzr2Pq�^c�Zf�?����Y���7|�ݩ�/����
�mk�S�þ��}!Q�*of�e�?�P@��~C�E�tۡu��E6�;	�k!j���8�ߧ���Q�g[|��!(�ZA�������s�,�w6��& ������Q����iBޗ?���~<˼��Aq� EV}0�
.�[��<���y$y��Ǿ:�#0(���� ����x�L �l~,4���?�B�bp�N���8@1���-u���5C��/0z^$O�T^�nL�o����n���E(E�����!��	���S/����}l��H���ն�☒�Η�R�N�a�WK�܁���?7�}������#����d&S�)?�,^;�0��#iC��}Y��uI/�efrF���N�NK�R7Y�l����Y^w��@����CQDm� K�6=(>[[�V��y�nӒ�h+�_�8��Ugh$�;��r � ����]9���n�����'[�_��|��U�9z1�V.�$r8p1@z��{���f�E�R��+����;�����\��lV���FxQvpH���P�V(�X��B*cGk!JW:NOU�
-�����n��?���l��Zv�R�E��%:N� �G�>�[�N������O222��b�q����
�X��ܪ�R�?��Y�
�O�ex�Q���^�3Í��\��텼��oSi�ؘ3+��)#f|�\���ڇ��,3����ղ�QbT#��@������N����AV\ύ�����Qdvf`�7�33�`7w�f�~��`���"ٳ#zE�o#�Edp��n����i师.՛�,��yu���0w��/1EhH�'�MU{B�(�<#>=w��N=����^}w	Xj��)�m�!�f�7g��~�u3�U���gY"}���U !�Tmo�>�^�{�G"ܔ鹲�p���	Q�7��I8�R�G��\��NͿ����\������"��ÿjh�ѕ��rH���vԶN!,v��������A��
��9)���.$��@h3G?AO�����2̗9[)S��c;�{!���B0,D��$���w��-�<p���`��`?�`�Mr� ҴA(G�[G�f��i��Q�vE�N��&ť�ϝSߟ{�JU6�I<� ,�Q{ɢ�,��!"̍lZX�T���ݵ�j$nVD��dLT��10e�뢐ب�pī0��_��ȳ�4���fs��&�قT��dҊ��w �G���8Hf��:�A��7sK{�F �	Ʒ�WF��M\K�Qw)A�[qB&:���v�_ld�/��Ǝ'�x�� ���u����C^ڶ(-�� rW7�r;��S��G;�#�B����DDD]��J5WaL1�cT6Z���(=M祒�e���O�cwW��P��?���q����?/�����-�����V/�fcSȊl�逩����S>�����S0�V�� +���`�q#h��o���/06��خ~�l��4H":�@x�T��K�Ѐ����ג�f� ����f�0M�}	�,nٟ�PЏ��(�����X��o�p7ѧ�P����l8�a�x1�J,���v��	�=X��Ђv��L��)����p�KFFb|�F�$���a�j�;��I�9�!qC�\۸�Qs�	[]���3�u��s�Wy��3�|���2�����s�TO�U5)���,��E��<K� �Aؕ?�&���Bq���.
pP��� ���܌>>��B�M�AE�=]�����5�
�vFʘ'ˌ��oO���¢�<�WH�VOFU��D
�
��j��\�u�Ӻ����yk1vRABj�����m��:i��2�`��j���dz_�ت��ֹ����3���ߦ|��:�r��Zcqq�)�n���?!V��M���{J(}ӭ4e�5��m�Jղ+&�,�0`H���/者<7��Z�}�0)Qۋ=���+Uc�����n>�#�6�_�tD<ś3S��#z��2�p�c��·���ד ��I9g���+���a�J�Ah���D3�7_RJ�lgJރ�S7mo�EUII�_q��
���Օ3#c@�Z��]�/b+/<�4i�X̢XSo��h�k�'�*7�Dȣ2�oZ~g���:���&��1�x��j���b���h��%�g� �5��K~[�K�G?��_KI�۬��UQ�^M�fO����f6S�&�]$��C3a�Y��{榛�}2�Eo�M0��=�a�[R:� ��dT/������l���;_?�"-�jN2��������E*l�CJF&�m-���K�Q�0ѫ�3�æ��#�TUUS��e�,~�9������x��#N���봨D/켅�|웜������&6܈��
�ML�G���>�і����T�>�Fq�z؛*ӂ�΅�K�#c}���TaOT���m��K57��$���̛���t���&��y���܁9䚨��ihW�̢���b��~����!s���I�Pr�uj���<�U��g�V�#�D��w�T��=�Vu�GC =P��pbLY3��h��,S���#lT{J,�X��%�����Ma҄�-ɖ�Ӧ+�+3��|�$՟����M�B�Exi��}4*#���d`�ZUr񦣤bs����馘�� ����K^n�����-ڈ�A �S�.���I2�3(�����loۯ��g}�.���NP׿�Y�"�����84�w�o0�"/�j���$���&���-$ue��67=���0���Wg6���e��|p�5�a�p_>f&�Wh�R,UM�X�f�cM'Erp��F��am�Г��A�XiqsíF���Ja<T��p|�T��fC]�~wU?aͮO��l����z�*���%j��hF�>~����ى,q���+��Ϗ��a�gXCf3�!�/��e~9�Dr��ˊ�D���J���M.�p�V�������α��(���3�1I�3�h�1�K]CC��3�ml��뛚���������*1C�T��s�q=�r��Ih�c� ivf����~�B����gl^�]pj*���Č��ۼ?Z�T�W��1�׽|��5��W]_Wq��������Ō����X �:<��˛*a�ozL��L�_2��fL�+ھ�Vv3f �yByjj�2+�錴:FΚ��t���|�}TXs���kǤۨ��<pf�[[0i#�/�P�8����|��o�\����Km919򨃮����-]���� 0�i<	��!yV���E-�/�H �����`�M��
�1��r��C�:q�mV����2�4QO�tś�v�\o��L���]肂.
�Iw��*�	K��S�ݒ�\jR������4��c�mK��K��>����$tY\z�jl��uX/�-HW��u���z(eнѾ�${�� z4+���II�@O�yt�GCdf�f�����º'�V��.$��w1]p��k��h/!���.C7�m��J�FO��^���G2�	�	�#�x����"�M����%+#�'���r���e�=7Vu�2B�4+�y���|�F-�X�E�"��B��d6E-�y�����u��F[�8 h{��7�~�J���E�P��sr�(��"�X6����bw��= ��F.�`���	/��[9���J����[tt�-������}w��B���li����,�ͥ�E��=��5�>Y�nM�X6��C��\B�D�udL�&�D�)F2_�-+d�����-��	<`Nm�ǲ���%8��2�;vgׯ./�g��xy��-)�d��q�{E�A��}-|b5y[�����CG��pi�rh�T�$96$N�@1�ⷚt8G�w㣢e3mWo2�+�/I0ȣʲ��̳=qmmm�k��+��S����z�	!��i\Ɨ��O�4�)"��&����-&
=�8�����(�5�)�o�X�b.T:��i��(C@��ՙ���u�E�Em�4�m���a��T�:<�܊��4�b���b�JJ:q&�E�F"	b�v�+U���J7o�:�|Ӓf��뭡�̈́���B�mY�[.�ށR[��'�Ч+ ��ɠ�Aɵ�~�\ta��H'7#��l*�Ŗ��
�� ���ύ�O~��Jc��vT.]&����M������o�FO�D�e��ߛ6��=�u�[~��=(	���-ӡ^�vm*Y��\ڟ\�i5�����'S��܆aooo,~�C>@ �}�øV�I:]y�f�1'�RrہֳO�p/d5+T���s��r����c��L��k��|o�I2��A���4wr����f��7?�ё���	�O������̜�֓?��;�M\g��a���ō�WhGL�(��I�Z�9�x��[~�vE2����O	U�B�� '��ٶ�ːP�֘�Y�?7y��r�(�ڻǬZQ"/\���?�h�Uk%�ufdf���A���A�ma��j���Aј�8]��z����~wz�O�M�!�w��o�	���"**(�&��:&��%7wp���l�����440"u�������0C��*.��B���ƥ��D�<lh�I��;U���ҋ�Zo/o��A@�Z	��G/�Y�ɞ����-���]��-7�U4g��b����/�5c��:�D�Q?)۸���oB��c�K�����$����	æ����D} &�x���6��3��v��_lҁu9H���B})����]1��©au��}:C��&�&�e��$ųM�'&'��L�ց��V�b��oqA�f;���0S�t,s������韛���VC�����:@����7�|��|�u�/Q`$�X��R.t��b�w�D�T�V��+E�*[�G/̚ϣ 9����sٙ������6E��`yl�u��S��}��D�_dE2??<���<:0Ak�#�����1_:GA:^��d�������N}s�ˋ'�ty5����0cb��`��Ľ�:N2Z</�zrv��E��㱔�	����Q�v�y��ďV��Ź�c�R�pq�\t��v�eMK"Xa�|�� lެ7��d%��wT#�CrֲG1b�8�`�����-�ջ�1�5Ir3�������f�SՅ�$�7y�	dC��f�Z/���m=n)�L���;���r�>v�����f*�g>��C�R�W*7��H`+��n��b�
��b�E����\w�����i]8���+L�i(4�T,<6�T��8,vrwg��y�)��qP��y��GG�]\�ĩ��o�./��D΅O �������St�y_����7���-$1[��H�-@]e�c�ߏ�^L2?���!7:\�S�h�Cj�mx�3Ĩf���q-��R;�f͙*�:UB�}[��gm��e�4t+�WX^��	��>0˩c��fJ-F��my�l�!M�脬22u<�z��3y0���?111�U݂%����E����/b�s�6�(h�ȼ�҇�r��p-z�+?DJR���`�0��P���Pc-��zjVf;ǹ�}�ޤ����W���i��ߨ��up0�(�[�K���dJ�Ƒ�*���)�]��D��툹���͘f3hD��̆���P�p�Z�x^���Y'!
B���n-Q���4B@��^�NՅה��"_~�������F=�������8�M���Z
񯕕�	�zz}�~��<�l��q1KR�J���z�;�Z b�C��:Uc]c���)B�:�Q[�i@<�����Qsf��꘻��;w�vn4|�M��Lu�<��3�^v�go��B2C<L���`�;���c��Pj'�8�����%��S�-������D�t��6�������֏W@B���s)()}������Z��5�C��7�^d-����'�L��Qe�9E��d�P����N��ݽ��d8a��q=�강͏�:p�ϩ=n��B�x�������-I�4����x)f}0�@�U��oTC��y�r0;���x&2��.�Y����f|��g��S�χ�#�m�ޠ֗�r����iKE>ߓw�������آH��s����c�ڪ������N�a����e6����9�����G�Un-��(1"�p��snS�x;w�2�U8�6�}��޻�f����vo�f�y�Z0ڥ�Ѷe*j���f��Խ3�B_�����{<=\Ac�J�p�"v�Ј`C�Hu��$�+>���fs6�N��.��m>sپO�w�[JI�'������!1qW:�MKh����BU��ƣ���O�^,�'s��_?V"���X��6K��M��G��l�I�!1 >M�����p�pꏹ9�ǋ��9�%"Y���c�_���d�}[۷j�VaL�t��L�.cm�Z�Z��Q������]h����_%��^�����ۤ�QUU�S�� $������q�ۻ;��A@��}%�A1�iA�<rX�oqJ)�]�V*Y�L�ܷ�_ǁ�W��+v�_)1!���F�K*�?5-��"�[,*�K���FG��Q�ՠ��2����E�ϒ������܅W&����ִ���m\������ￆ��5��Z�"���Ͱt^j�_h������a����6��ʣ�O��JK��,G��Xg,08z�G���:RU?d�	n=�L�Z���!S|��ZC��!�ښ�w��
����D��֨��κ�Yڋ��ۓص�Eiq�G��X��pv��I*}ܽM�Z�rh�WFU�f(N�\r��:�c���8ߜ�>�X�g^� ��_����h)r��f��i �i�yt}��l2�ܪ�̹�B����դTѱ�u� ��J	.��� cLA�H7�M��B��嵉�IQ=a�nr��,�H$^D6�.�	��Pf��h�y������z=�:w��S;�w�~,N䱉�^_AQ1}D޷8D�þ�60,S�4��~���R^!E%� _���C�7��o�ܤ�b�Wq�����U^� Y �,�ￖ�9]��
�A�˧�@O ��D�&r��9����p��;���n������X\��8����@��燐N��=��@�zďZ�J�[�A|n�HN\���@��8���I,>O���vJ&Z�X�I��=��7/�(9��'o�gN�׍%�Q�G�_]���uT�~|�'���Ϗ\^^��bv6�勛��w����HiY��J���*��PAK aA	�cJ�����(�� �$���2$�/�`H�緵���L�X~=�	���; ����ē�c�8.+_���9�G�&[ȣ�S�h���m��׋�x)�����.��UN<o`p�LZ96	oD���̜�;��{u����v�.UI�!v9�A�����D�,7x\�Y��2� ���f3[�ǪD�{x����_�����>#����/A\�����.���O �"E/��ˍ���*�W_{�GT���f(�������:cJ<��֪e+$�,�ZD��.�Ӊ�Nz�qq����0����%;c<�O-@�~e�c���=���A�]Ψ9��M�n���{e��p�&7�����>��U����~�j����%z��].=;۬�L�*AԾ�s2S�����~��9�awʉ?G��"??'��ѷ��X�]�-���_A��o3��W�.e)		��W|kC&���m���f��xr>]|Xă��=��2ŬO���+ǰ�L�RT-�e����	��lN�e<q�SSS{���e����
s�����7�L�jtt���.�;d�7U�U���}}$	�G�+��2�K�['r3b9�o�Æ�v=?�AG��]�+_Z�wAإJ@!�>�@�|�y���?S�9���L�s/%]ќH�B�-���"��0�\�t�h�%�'xb�_�j\����~Kl���:Jء�n����b���ڻ�?����~ ���;�d@�O�5�D��Ӊ��b��H��N����?:��Q��(J���0��LU���S� 
��=ٹSd��qJճZe2
xQ O�A]���v�M�)\C��G8$<��Ǻ~V..���Ο�C�LU�nTs3��b��F	�b/�yq0��Zfg���y�m)�EQ�Pޓ�I#��H ��V����\�ƈ�����v\ ���np�����ˮ7O܄���kik�QMOO�R���]�ʲ���w9 M�a����w��������3Rѧ����a�<��@��G���R>v�$1�+���g�^�]�D���S��}��
��(�\��Q�������&i���O8 §N.ܝ�V�zl�]E�Lx?S!-:y�.��P�9���(�G3�=.1ymaȂ2QQ�̄��>���!���rڪ]��W���BΒ?HѶB/*�h�!i��"�Яy��FSW������24���%u�#IC�\������I/vp��T�p��-���}A���soh�'�ӗ���_��59������z#�[�P���1�y�)��^a�=ӯ�v�G�ѐ�:���yP���i�b��{��ə7 ޘ(U ����;��ݢ��$���m���p���OSN��Dm!M8ddc���]�#i��c�[��aW����f*���r܋\{�O���SUK#��&G��9G�	080/�R��0�vpAEy�B�3l������Pu��/���WS�+�ej��]�`Q\�X*֊�	0B侇�s��L��s-����,������ /M~w�>�^��i��ݕ��t9 M�de�]T[XXp P}S��	٠��r���G��O	cd;��&7�г� �7и�(�u�_ʌ�v��ĳ�fnm��n�H��.�<宒��L~��;��������A�'\�W冭n/�7�$ဨ�񃀑 3Y�=�*Afe�>T�+�����bx<�s��ȶ����HICt�r��� �\|�kb3|ťh��m\�����WXI��
�.A�A�K��1��j:�Ԩ^Y<!R�*�C[�S�4ih�6��@��|�܀L��}bUz���!c�W���I[\�V��M�K�j�|�h�oA�>�L�����)靁 �Sc ���#�>����2y�3�;/�;�v&�]��)^ZڅMW���I��<~{2�i��,ysU�1�+� =��v���QG`�ķTu�G6��uf�b�@�M>��Y�2�疵�3��A���J�Gq$��YS�]�j�]��J5h ^��d���\Cp��)Ň�E���.�@	��%|r�l1&�N��Ï�B-�?J�.�m4-ol$â�3R�q��{Ϥv:m�����b�,�mX����\�PA I��K�d��`�%޸�U��6�`������F�쫵��n#Z�#���|tZ�BS�S�T��Z�l�}F���׮�dac�s+��o~��z�5�j�L�A������?�,��rkl0ᾙ�OʢQt�p4���۫&"_pƘ>�atlYE��Fg���Fլ����,|���\h�S���fI��k\W�����/�7��P�N�)��`p�����0ɂ�lB�U\m��������ؘ�+�p�>_��9�)��	�K��)A��(��d��_ul0ZR�K�X����7'I1��Dk�S�zK�?.�V��9;t
}3�<Dk��*��t�J($��X��%'*���m$
�N����.@|w�b^ �omi�����s1T&����y���3�!��I^n�0k\�uX���`:??7m�䒣s�����G�J���E�0T�5�J��nRM�w��8�����������ձ\��i��U���Ao/����JIF5�-B����.��q�zÂ����%ݺ����ِ�t a�ĩL�o��o���� _�½!��2)��������᎒�(�vL)���Gi���r�[�������������������������	���6Ϸ:::�K�l�Th��Ri�Ir����bœ��1�����Qs]�Y�8%���<�߰���qPJ�(%9u^��y��\y��S1�)�'Ա�8��q�}�r��$�L ?= ���T#ן�J�<D9l)	H�i�oArf��t�\�K���
��X'����~gN����f�vT�������͝WZ*��*)O#�3ʻ�7�G��ZDD��Ieǅ�`���6~�<`K������L��N2�hs�I�?������	}�&���1F�u�t�(��B�x��0���J��r��0�,���K�K�.�������|�ikm����ؐ݌/�
��%�6�]��kE�4�Mn5"�Q��;x�(�pVT����"����p��j.�ـ�I\����E��L��F�k��o0WO^>��F�H^��#y��cj�c;:==���Y����\���l�w~�%'?���E�FEú4D�I�w��Z�/.�,9�$�+M��ҁ S<A-�Oq-�1���(
Ó��T�@�	����#/���Dc0��S�����uGlׅx�B�xm`�'��O�-zP����H���^O�A��g�j�,�Ᾱ�y�q��_t6�u?�������/ZX/)�|��]·܌��㝚o0�*x�85[MB��	C��5t}�}�^��E���C��R�����gx��۔�S$�vke��U�pÜiH�/�p��滴	gW\շ�d�t�Jqr�|����C�8�ˢ�{�+��9�Avm��ܼ����R蓉�h��]t���w�G��V������ �#YF�C�}��շ�9?t��m�p�u����)���ȱ�}��?�ތ��Ye1N�����t��r����Ȉ��ac1$�nD�C������n�dp��}@o�ˀ�3bi�l�f�:�O�'�[�Q#l�Y)��3��Z����fU�=��c�v9�M9�c��3G�)��n�� ���GIR]���C���Ӄq&��5,ދi����nh�0f��ix�F�M�lɕ__���>�rI죲�z�Df�%W��Y�퍩�@ <rMK~@>9yh>3&g��̓_�v������G� ��K�,<|;䀒]�{|�k&B ~�
Md0[��_�_O+h0�L̹�� ߅c�+���p���c��Z�}Me�⃛@�O0�3�~��4�C,�׿�䦶���c����]�~!@�3NK�X���J��)�_	y�!)��Ī1��W~���/Ȟ� ����V���j/0w�������*g�]�:��!�'�g�f
D�O��@)~������ҙ\Z�U�Y����Y8&���U7���@+*x�ٵ��
Zp��v=n�������z��\���Qe�^��j�FFF��M�� ���Us6M���ʚ�i�Ӹc|���63��s?t�|}|W�.#�sێ?���)k�..8G���X�G�c�[�{��v|���������F)"B���ji9��*�R�^�i�D��f3��KȮ��MMMʹ�%d`p�`D~@�|(s��+s�tY�!U�SK�,	�JB.M�^�1/\ɲI(V����d��:Æ��ga�pʭ���xm>@"UU9x�
��lTҧ���@ Z����066��v!{sjEW���������/������5սXRr�F)+; ���m���o+�t3��J�b ������H��0|��ȓ�R`b�0j.?{��^RQ1��L9��/�u���!��駵	ؤ�pl{&�[A�ӟd��JM��z����{��f�-�/��6&���5�=l\��>�ᑭ�k׌CLl��ğ�_:�k`@�vA- �������N(XvD6-��?�&v�+����G{Ͻ������,�w��KN���nnnK+�@���zWW�l��v�8��Xh�uh]�*�2�"qܙ�LNI1�727G�k�&u�2���jY��!���)hS���߮,�%��p%��J�:�;��������R�κ�hV�v�1�1�ې{��`��7-�Q�R�a.)���)-m���w��ܔ-��]��>[JTmd"���[&��ʊ��̻��.�bE�k�#��0�#���8�����U�X`9�7U�E������f�I:��~�Yޒ�lb�iT���T�%W��]t=q%��ף]��$e��E�rL��ih����d���}*I��[]]�,b����j__S���7��}��'y�Ғ�䗕Y����O	�G�jz/0h�Kݢ�w�n&�l;M��~���[�8�[�f��ʋ�#�ذ�?�xy%w4�t>��A�*���� a����'|ԲϚ�l�;�-�_�F�s��f�R�P-��-%�7d	�̈́�Bƙ�(i!�;I��="��m��8и6��(�h@s�`EV�"+���)��mg���p%�k��r*}���
�J���;<䆛�i�M� ��~��O"ek�{�4����qQ���
s0�(ÞF0�A---�1�\i��{MY?EC�b��ݾ�?����3痗t�ud�S+��}j���\h0��>�����_6�C�໿�1<u&$$, #�P�����ֶ_�wQ�{t���X~I��qi���, �#��;�I1��}��y*!4n�0Ѯ\����ͯ��&*���PC�goo���頦��S7ڴ,i))�O\��@���Ҳ`�.�$F����띹�����{��dzlC�_��s�&.����Mq�jCb���	�\[�"�9�R���ӵ��&���2W/ߡ5'mr(( ;��K,��y{��g�cm��6;����)L3��~���k{^��E;��J2T�#��Կ`H�$"�^��vGp��ow
V�F��1�j���_���nT)o��3 �'w��C?��].��	p:���+z�������3�#��������"�	�i��v� ݠ���s-�:�sq_�L3T:{C���_m��3TӶ��40����6�� \@d$��{~Gy&���C��{Se��4O%����#�?�`��}��f*f�!:I�Z�}���鸊�摑��<ZT��G@ �6;��2?��i�M��kl\%�X>6d�l���t�8"+ЩjX��/ �V�)�\��q�o�o&{Δ��h��N����_v��<?���׿�i�<�M6�;���;�\NX��_��PٳZ�[��hJ�M�e�¦
7�;�2vh흰#�L�K8tJJ�]M0�{���Od���u���e����dƄquqYI�ȑݿa&@ H�OL[~>�B���o��B�!��8��e����h�J���)�N��K�灶���StT4���:��aj��9!��*�6�{	Aw�32H`D_c���9��:���j\�l:5W����(�N��n��qGGG�����+�B�b{' g��3��a��#�^�B�����@��o>�ЃζF�*�x2�xE����=�#�����x} ơY��,���uV|��	嵔
���6�NA��N�?�gy�������i� ξ0���eA�v�����W�O��/xQV��A���>"�=p:��
	��y�)?�(ι鮭��C����!����3�~�X����֯���רڽD&R3�hMI��>�»�y��v�o�9�V'�ҔeD�|���4�&K���3�l>�nGwG?��ĸHa�� �O�� ��־7B�s"�1�,R�"�G�77��F�B>���4�����fx��� I���&w����`�_k�gj�۽�tFPPw���`��Ǐ��_���|}}��)�����o���>�V��3�Q����.�?U���q�R99�Ţ�M�6�%P�n�+����,--�N��![�N�?�ᶺ�t>��񅆅�` ��ͨ��{��i�{PaЦgsɡȎ����z#�&+e�L�ˤ��F����۱���ܥ���_���8��J͈��+�6�����O�����un���G;���<���0�)��U'ſ�"���n,�xA�h���P$�i����b�SC�]d���V��qP$��9l�;Ƞ�Iæ?��O��p����rr%�������^a�t��BGZ�N��^��L��f:.��e���0��L%lC�J@1�Vj��Nuai�Z^n��܎w�!���Κ�?0Z�u�@�.���.���g!R�3Qǝ�Ke:,��5^:��$��(�Q��F؆O�3����l]G��oyV�[ZH�� nN�`-��\lu/���'�f�I���Z����������N�7}���B��R)��s�t��#��v]b����N,?�����c�:�g0�%0��Gb�u�п�ͭ~��ը�L�S9C|���pv��Q}\�\Pw��]`A�wS48�giJ:M�b'�N_#�׷ۂ�1��L��U���� ���g�u�Lf���Ps�#C���n�BLlƙ��[��P��g�zs&��z�Y�[#�H���B*ŨF��Q�|�c;We�r���DO�Cy��x3H#+������AЎTT\L)�t�5Hԛʢ�0��8��<)�`���Z=:Y\RR0���jR�� ��ړ�U����Z�sK��`�x�!Z��ëI�Sv�uz��rp���J0�X�W���WVQ���� �-̆SPZ�V^^�Ns�1�l` ��O�*A
�M��b�}�ƈ�^�����ӏ�Ŀ&J�䇼
/�E�L%@Ps��4~VBP�pu�����3���Rl��u���]���r��0E?�m�JǑc%4mo�r�}3��^��e�A�[�E�+��W�#̼����J�d~�k��/��������H�X� P=r s0�yUU�ִ)������ɨ	��9wT����]GHII)�&�y=AE�!�ٚ/'�"d�P�[��n���vZ�0�0]�)^e��}�hAA�5tY^����1�wU�����ZX�pq�����|�k;�*ho�����fNV|4�T	��B'��ZS<`�u�Q�x�t�&�+�4ц�x\#��/����^��zкR�d^s3ߪ�����3G���,�Zr"$(d����xe����5���^�݊S3n���Am+&�[sM�19"�}�� �!���e�/�C���Zx�/����М��ta܇1��{������ �CCyH����;lH8-2q��u��
���[m)]b�)���Q����M ���#P2�#Q�wك68��D�ϥ���*	���_C�д���[j �y_WW�5/�x�@dR��b��� �}_y�R�OG8=tt,LL����כ����I���p$���i�a#���P^!���Ғ� ��_�2��`^�А&�-f�ｽ.��+筕�T��-MbM�L���KY[3�2w�H�A�ϕf'ҫ;�� ��M��l�wo ����o}�Z�X�G�tv
z���H��ʀ�O4�h��T�� ҌG%�r*c�ܼ��RRRo��GG�Vj\�z�ׇ`n�6�n�`�k����, h[T�xlqNk��g�����{�4���!wB��y�!�0R~�Fy�}@`(q��G���3A�lNK�����Lhh��g}�đ_�S�11��?WR5�i=??�,WD�:�uO9��;��D��a��:�̹H�O��!��H�b`��H��(�@lu�Ȳ꛷�kk�K���ͻy:�ㆇe�45-�[�9���޼��g��q��r�.����������$����w�W�<�_�*��
ev�0����b�'��� e<�[��w�ᠷu���`@����@����\baV�lmYܠ�R3�%��#ha��ֺ/�������	^�G!��	Y�l����D�;~�_�i��\�#���� ��qeM�q�Ր-�K��ph�>�T���v��p"D�����e���}1�*zm59�@X [��AS(Xm���J���*�.��tl��]�5�n;͗x��y	Ŀ<`l��#�e) G;�2!=8�D�0�8ർ����q�ߎ�p^�R:�T�����d�x���h�kE:pa���L��q��� ~z���D��'*�?��ħ'CJ;s�O����َ�ڈ�J�m5�I\~�k����Y�&�<�q����VT�,
�h���[�Ǝ�!��ss��\o[��u.����2�һ�P2��ޜ%�7!�+ �����GW�KjqM��6A��^o�|)Y`m�i
�a�L����V�M�0 i������X��{�0�K M�LsqEN��l?�9y�����n&wn[�@��
�wKa �������V��O#��\���4�leV;������<�D�����y�F�[6QYS3���q�>
V>l�C�N�����Q��Dr��i��7yqԂoë�;�����z,,,��a����l�g�^%� ����GG��z7�J�����r�/H5��QM0�Zɀ駪�:�!�;�708�D��4^�,�K�J�i>���J����+ʹ�3��3��KM.�������hZ�0��/Y���zvzG���Hچ����ԟHql'>���ڒ���^^^�a�ܳJ�����ӗR*������zuQ'�W|�3�wU&:_�%^����|�vT��.�;m ��a��_��er)g�nnnZ�ۇ-�rv����e��l"���m��^ER��(�$�(���jG���hY�Tn8��B7�w��]z����Λ��t,@����Ay��·i3k�ɟg�Э�f�~ �e�d��,Qy���.�e���n�Ly0@��]��:�Ȫ�:%.Z`��t��&щ3M/(�b���1��;)����E�d�D��e��F�V��{`~�̈��G��f��s���_�*#�q�n�m/����lbܦ�iAT��y~yG\��]R���\���5� �;�ٿ�o��� :�fhiҰWf��K�vvf�ZP�kb8��vH>�]��0��4l��-=�HNM��T�<K��p�3��i7�S��1~�w�[��`�cx�0��"��>C���-��U����QM|���4�WB��~I"gM�;��n\�S�~����
�8�����m��\��C� !H������-x���{��5����������֚E��g���ޟTUW�����-;44PSS3q0�t��:jv�Ò����r�1؆���I�oi3��Ʋ !�Z�2"8��>hll,hg�����p���G�����Z�AQ����Ϸ�T<8��}�P�1=��&(x��r�{�u�MC�>Q���)����XYm}�e��״��`� ����l=�H��m�7{��_bp��C�A��x� �tS�׍b?r��5V���-�Z_(�Z#�}�5��9�$M��h>�+�L�)yN]���l~$�YmT��T��+հ1?@p��
o�g��M�
O���|������s������QdT���~����ݐ�g�=BL�.�~}�C�Ռͫ��0Ǡ̌�͕����rK3�66J� �
��cM\�Q�,G�oH>Ȑ#���#e�D��̬ۨ���@�Ȅ�q=�5P�!�)�p���8�;�6�k�!�oM���r��$54p���S|�ڛ�����f�SH1�:D{ �[�t��Y��u���Q�e����c�����vij+�Cc�wT>�bi�VZ*5}��;�C�RI�!S���_,��𚆧��4�@��UȠ�����*�l E:ͯ�aŃ�u��ʴ`�蠸���m���ƒj�����qg͉���0"�g%�S��?E�ި�2i!��Tٮ
/9��~��S��ښ��8�Dc�_4�w�E�4�A��+ǃ�g�ப�an�;�L�$��d��r����+H/֢m�.'�$��	dn��ݽ������v�����XT �P�A�r��}�֯ϴ
bk��*���*GT� E��ߐ�~5�i?O��������r�0c�tȞ/@<�RR���0O�9}�����|��#J�ғ�+�TP+�z���)M>���T�}���#i����_s$��Z�i �d�uT7�-E &�m?�"�V����(�?<�~�|��mp�%<�^��^x'� c�C�|KY����>&
B��Lq�Kʤ����#�/�����Y�9�4Quuu�22T�G
�߾��5Z\L��@;�m���-��I�+""�$*��B z��Lq`���냺�7����&�2O?�p����L����o%I�:I��Â�"�Gl{�+3��i��CzPQQ�u�E����*Z����&���Ĝ�8����\/G�'�0{�����y͔�D��a�	���T��}������_����a��<����H37 Juk��.gזe�ۻس�+ͪ4!4v�PǸ3������.T5ӟ\会,	���v�V	�rܯlǦ�������h�G�ϳE*5_.���Z����� ��u��hB��3���?� ��k5����*��?d����L�Ĉ��Wu�S̻�>(�/=T�pM���T ��\^��j��{��Nvmj~K��~���~b[]��ݰ�#�����fN\���I�6a%���UQ��k�ֲ �j�o~�{߄����1�ɫ$J	�%vy�J���i2�tu�QT�������o�]7�uv���s�r���gl�������]�����xb�珨���:�ٝO3<~z$^a�Rmil�n�1�Ǚ�u�c�e"-m�G���	�⧻�l��U�5s}�fk�9�� ��~�8�����Si��F577�D�Y�	�߽�0�덭*��t��_�*����S��C5���bRܥ0!���Fi<:���9�����+�1��2��͢dj|��)ͤf���l�f Gd��r�>����L�F��'o~g�=[�c�I���!�zx���п��^[_'����XxHϵ����2���ľo���ZҺ����m߿O��Rݾ�c̺\U�вg�����|jHf� ���ed*�ǺjQ]���'�q*��`��RQ�#d����p���#��# ��ZZ����muF9��P4���YX�MLh�N��u�YYY��_o4�لS&E�^)p0�l����N�ò��8��S�kd��d��}{���쵁���*�u���F���Ʃ�;2�#`B?7w
N���QS	))8@#:R���|i�Q��o�|�)�O�~u�_Ad�x'��`�r�Ntr"lY��L�(7@�b�"Rh})�C���FDn,����ov��w�|p�ܲ�.:��?�"9��a!5��=�������<����U�o���m�M&�zeee*0���,�,��]ʊ�xQ�#���Br�x�_罦f�,uB������R���G���='CCCʽ��l���H;��!�4 ?W{佉;T����>�l�m����Bmm�ݖ
��Q�Jݽn����ۊ{ɮ�o=�� �O�Q��u��6$�v���o���xI~,EҺ�Cv�\^�njj
Z��<�Wڽy�����5?�U�� ��yF�膑V�;��\�Y����7^����~qt����kY�Oՙ���+H���"Z�`H�2�MHL� ��楖X��*��5a���Y�0L@�c��.�YP�x����\�D�֯��|F��|�(�U9�o�f]R�pg-�M�~ �1��!PYl�������}°kj���� ��ų+I�`L�8��C�5��f���c��t����g@(��ңM/���uI�������R��H ����M2Nv��}�ڌƧ��ϣ���ʫ�@����"}������2���ީ
i�´�a|�=�Z� 9���oafX9d��LI,����f;�K�����ǛM���*{q�9 =���xnoh�s����QS���D¢�"zF��R���H�U�iEm\���O��G?f됿;���$�xY��b~O:i�AG���|ú��{���4�x�Ȼ��q��U�0.A��Nm���}}}��=sɟsé� ena� HU�������}�i�يͱ�l��>�9-н��3�B��w��+	�eb(�{XuA\�v�92��3�0�~Jɢof�t���Y�v<����	�Z��sm1�qT����eͥ��l�(.���ێ�����n��*���T;�b�''gѹ��+�f�gƷ��.��}�frb�GYU5�ʌwO�]����z1*<..�+����o޼�������l%Ad ��Ʃ�U��c�F?��@��}�=���W��|�5=a#�����91�����V�J^r[W�����Mdi=A����'" +����f``���� ��j���x.�V���*���>G���A���{l�X��nǔ�qV�c�t�3|i�S�w<�S��-C�ܲm$G�������5׮�!9�6=�$��:��.}Quu���2LTxv!�h 3�&�L��p21IjiB�i�0K�ަ����/�jO8���R�{�� }����-�e�BS����°�$q3v�BEJ����C݌)α�;Y@:�tGRM�`��p����y�s�5(&�%(urZ�qd�/5�" ���h+�Ã8ν�=��B}�L��8��<	�m���B�wz��f��pr�в��@��[��͛���n 9]\��b���C7d?�83/���E���׸�[.�l���������5)�otD�a%���G�)֪�5�PLY������䉺�k���A ^^]���S�}*����g`��ma��	�2*&@oCu���9������X�\\���u���� �Е�K��������'q۟M��[�� �J鈙{`�؞�|�eP�~�!`�{j&$�B>������ 7��*V�|����^�e�1Z	��d@)�B*�
7�z�ܪΙ9
�Y, ����cb�++1"�{�[U��*���P%��Qi�[���7`4��9���<���F���5���똣}K#C�M��v Ͳ&7j���fc༿�l�?]�="��9Ʃw��pjՔ��Rn�,���:+�=o��OmװҹȶM'�Rb��'�)�IZ#ү�6��;�b�蝦;�؁'Qi�Ln���^�n�x�J � )���X�85А�����~{�:�ħvP�*g��>�p�&q�jz�t��Q�r�54���+�3��tY�@)1;mv��ۑ�9���%%�||��})(*~w{%�*ή�}�\l���͏�V||H�����oSY(H��|��M�=��]���z�v���RfP���ņT*�"�qܷ�oqyݶ4:mU��z#������v��~����H(���[Ι����,�[/����;�a��u�*�w�ށ2GC��M�Ӂ�ZY�SPVfm���Yy|�`$;}�����#퐸�p� ��6��/���K��dr�f=���J��8�d0f�v�Fd�:��ߤ�yw�<��Z*���-��<����F���_)�����q�Cߨ��i�g�c �J�p���?I�,E��xc��Ν�"wHRb)�%�DSL�G(��9�h;��B�>����1��$�xxy?~�u�:���T`���ݥo]�i6!�~[�ef���)2$j6�W�����'?�"�����\�6 �q��:�|�Ց?���	�S���J21��ƒm��JpXR-�;|:|�DH��Q	�+��h2�omo��h~��؊��OY�����wL�%q+�E�լ�WM-Ä�o��ڛڡ�G���.��Mϓ��_6Cٞ%nCY}�ȟ'B'��k�s���I���Cy��٘��ʇ�@k�+\�ͳΝ������
LD�R� ��
IQ�M:�{{b���溿z��^HCD�`�]h��ma9�e�E�Zd"��:����Q;$	�?�LW%�PN����'D/�u�ۦ�nf�AY�-u���\#+���b%)!��m�B�k&�!&�o\�b��g!���屍uSȶ�PJ�ׄ�āS{�jj8�P/eT�����<@w	�Zȵ��T�: ��.�z�s)�w/
��h�4HO@m]��%S.�2�s�UUU4�"bF�>{e=at�y�\��Q��~���q4vpy�>��J3!N�������nJ�&���⾾"�.-�c�Q���,e|$�=Wc/�tH��A� �+z��T�W���F�KMG��8s���Jt����2R�<=	��L�#Þ��؆� ��2�f�j�c~��`�{���ze}�j�Bz�v:n��k�}���s�wvv���p����9�WA%Ij.9�y�jl9K�62;*�^z���r�n��pἽ������IQ�X�����x�`#�[?��~�?�2K�s���d����`���ĶY�È���:۞���i/�6|ꋓ����Tj|������×] i �/)@ġ���z�P ƚY]NB���6�H_߽E^Mg����|oHw~� Bh�?1��p!)r���������&<)(#�g�gO�:��M-��^Cv%��m�U�_K�b_�����`A
%�C�X
yx��d1���uﻎ�F�ZY�ߏ��	ԧP�� j�M� �����v��W��A�<CD�ߐ�nl�w�tnsG6[�d�ʹWJ�i�Dx큁�����+�;l��^k4����������
c��d̫uҹ���#�ӑ��_Eo_��4�4H�NMM��ZLXk��/���ļǅ����eϥ��������ݣ#���i���?���~Ki���c���Q�H�㋀O��廪�~\�Ý���^�� <͸ �X�
$xcz*8�%@y�:a}�433#�y, ��p�"���nx�7��Bw��q��so�{�<?=�$�(f�= T��|�ř��������9�&Y�);?wz��?�#����u	�Ə��y�KHo��H��v���V��v�(֯y+8��lhk��~C�f��R��^>��FrQ6u�GM9����8۽������NTT5ZC���A�n�e�8��#Ԑ������!��x�{4
)}�	���R�!s[�Ĭ��0Y,B�rn���;���:��d�v��!cq=��Ǘ(������	j 	Cɕ�u�xvQH�M ��/]���DJ�+���C��e,���� FӘưj>W���n��6l�����G"���Y�T�lr>��4] 8��$�Т�����n�V!2X}s���8<�F3�&�lu�t�u2��@���}Ȇlk7����Ϭ�HCm����0Ʉ��ev2W�*9*ܳPv�Ug*.1�Ŕ.���5y'Hc�FP�gG&�r�=2ĥvg�R6�{�M�V��1Q}��ʢ��B ���͋�ӓ�l֏�]=-��D�"縋�T1��Pl$���C��[�*ZN��6[b��JrsN��>�M��ٵ���{ N�FxTl,k[;y�t�� U���Ⳣ�-ch�Wy'��LP�+_\��ZӤ�c�.%�ܜee��)Ťs�[��9@�f-�^kK$e�6�U?��G��&%`�������D��!��Ʃ�x&ͪq�D�W8��0c�v��f�r�r�Ѥ��~��v��T	;��&t�������Z�Z�e9�f+�49�u��H4���eZ�6j�5�.������Gpt��
oἏ��zB�[�W#roܞ�&��|NNN>�t�:�����J+�Å���۹�e�멹������)7ph��0�-gʴx�g�F���Z��"Q'B�8S�&�|mNC�v��#lrrR��6B�������N���`Շ+����6�L[��i�D�S:ߩR�_�#�4�j2�^���y���{B�@��'��/�kMz q�1t��	�u��竌f ���/���)5_nÊ#ɡ�_6��I����#"����ɸ���J�lƸ�浇��nI�X������{�%Y����K�d�����g�x�&f����.�v(~�e��4%���,�@vT����x��}]@^\����{r"�*N��aww.c":��|6po��}εu��� ([o�u"'��X}r8K�1��<u����~�:�]�|yd��M��g426��1��L�(�\��é���{����Q֝�Q�S��o����s�ٞYc1���@;5 _)S��WGZ �����W7�ϻNo��9��d�=��l]X�R 9�A�@�+�t*�R6#�s�sh:�%
�v#_��@=�ʓ�<^2HR�=HQbAV!�<�>2�S�s�o+��\���냀tC���1�fl.T�풄�hv`,�Ւ5� ]���?��7K�V�~��κxܷ����8�I�K���	LD�]�h]Q��=�-��=��˽���c�s/��KB��C���g���?4
J��c��"�o9vƂX�%�>�ޜ�'�=>������DKC~��A�a�0H4A����l���l���#=Qc1TGn��%���~cV�U^0�i����o��x&ͼ�{� ғ����t�Jғe;9U2����'��,x���	�`J8�xqmAR���NPKr��ײ���h}�Pbp��\�������*dGe9׫�'.����		}7�_0jXĊ��J��g[_7 ҹ��n5^.�͇u�9|A��X}�h�3�+f|]d�D4�ߙ���'��z��om;1���oH���X+��"����;U A+�u�%�����. �$w��-3�5�'(��=H3���^�R*�����
���f�:k�G���/j��d}ʾ�SA���y�����i ݠ�������#� \^]1{f'��Fw@�*N�w�~�KkZ�]w��p���@���C��C�a&>(_�����>7:�d���ȵ�@��^cK����K���,���;	��Y�W��$x�����9�����3o�F�Ԟ0U3�x
���9��&��k���F�2r��}(x��vJ�I@҂|_7�$�Y8��P�N��;�n�C@�n��L�\��m:�@݃�����&��ӓBH�Jr�7�$��l\\A���n�947�Dȧ��܂ܪ�����
FQ]�fEׯ�C�������IE߅i\�o<��*Q� 8��D��R�Ѷ1X�.�>��s��PbtK�[<�FU����@���.ϋO:��F�R�l�� �|�c��9H
�6��r3I�Q��*x� {����.v�jj��"c �����3�q�B����2h���s�n�#��P�!ЃU�FA��[=����[J\2�|+$�J��9{2*L:���B��O���B��KjC;�zρW���	ߓHזp`�>�!�Ѯ2���X泻W����u����R/�����7IO�ȯ��'ޖw��d��}{���G��8�6@��!TĢ��H$�~��S���sBb���l%�BJ�8rWjK��:�Q��pZE�� ��'��Ԏ���m���o��Q�r���ң(Hq@ۧ���%���C���$À���X]�0F0��D9�y�:p*��1��@�F���hq\`�!P1O��*�椠���Sj?��קp��xR]�/��i
�Bk�1�%����rTPV�����ϟ?)K/�Mn���:�>i��4t�!�wQj��O@���1~k��;��Q���y/�����&;3���gLx�!�P=!@�Q�QY.���ZX>�6��:o�N��AƖguH��M�ߠ��p��CyB�@~����Y�_�&�zr��۸'�;�}q舦��zt
�:�@�&1@�?����w���^�H?�!X�Q�p�'�-�+������p&\ �@|�ME�\Ջ0r��Eh���s5D�l����:VV�����Vip/��t��v7�r��y���	Z��74X�/'}��YW%�@r�
��0+��w_l�Z��O]��7a,��bH�$'p㓬��|�j"ݣ�$�7�̋�:�s���xxx &ym.��$$�rP�Gvm;t�9s�'��U�+�{5yNE��� �Tj��c���Pל�*\�1���� ��]>�<�k�t�yxV��k���_��`�����'�ߗvoۏ�|�@��-B��A(@��y����ls��l)�z׼F�[���&�I'����%S����?�A����fB�cBp�4�zF.0�Ho�]��/;:2GM�� ���2�&&���5�9�ʴ�V]�
a�����O}�R<]x���J/��ȴ���G{4J.���<!��;�{gvr�Y�ͱ��W����A'xs_�����Q��/���p#Ĩb%l��m:V��R���u�e���!<�?�&7��~T!S�Svٟ�z��R|P'����A�>�}��ˏؤ'#J��ʔ�K���]WnE8-����.h阾���2W�E-mF�V��Dè��d�rm[��x3#6�#H�X�P����0U{
S���%�f���)�z\J|�@�F��B�2����1z|\h��9N�R*k.- �!�#��a$2����s Y!�G{��2���t�rs�Wεx!x�uO����l�F�<Y�+Qb�m������N(D��춺+�a�y̲�����9j�f/)M�L���-%#)
��A�,)#��O�G�=e|�]ZQV#xB>�ǟP�Z�1���[��������:s#(3�^:� �����h�Ԏ�;�۲U��-�nD���UZ;_s��ŧ0帻�c���=_w�o���<�����sʘ����Oϙ9�Y�؉����K1ضs�>:%��X������d���5��٧�8]������@��8/���K�r<�����WN��y�����>���q����/u�M�JX����#bG���0"�ow�0#	X���c6����Z���,5���n��O�iF�y�@,��iӉ�V�!���w��$c�k��L�3K��c��t�ي�F66����k���|���}G �T��Q��"�7D"+�"�,6 R����U}?��q�����[��oé�l/�hWY@a�p�݇@�<\w�Y�"ԗ��*6���3���7
�;e�ڮb�m��0�7a�o;5NZ/�^�^���h�/À��(��<�8�~���4\��B�Bz\W�н�n9i_�(T�k:��hk״O:E����t=�~�	����	FZ����iNEh'�V;m�_��j�w�
�P^^�z���|���@�:��v�U��v�]ߥ�+Ъ%��b��	{�����9��<����nM<�}~�=�D�%%����e�0�%V�����Nkr[�G|�Y/۞w�B���7�����&�����(�T��8|OR�9��~UmM,C�U^����ol��mn��
V�n�d���*<�
�%J�h�)}��'f��{�� l���D�a��;�#��%7�~�ngj���vv����`������ͼ6%���*���s,$�v���-���ڸ��`|�=Я���o��]�l+�������>7%~�f�a��R�q)nl�����q-}�ef�����m^Œ_�4HP��	���^v]}b���/�[�-JB�"�{r��r]��c���Gf`<Ht뺅B۬\�C7s�B�AF��U����*Ha�cq���ܚ��'���ˍY������/	��U�vO`����x]s�[ܕ�D��r/��KK�9323�ݵ��H���^ƚtЁ� �K�[�9�G-�az�F(��2�/R8au,��g��>��u��n0��5^��	��h��ֳ�GM:��.G��g�й��,�E�~�����U��lSn	UKE$��I\P�g�e���+�s}x1��U��iで+�L�5g4T�n�G}R�ͤ��Ud*�r�~�߁2�����U.��XZ	�z>���Ru� yG�Ą/��#����ؽ�^tad����gi��[��ۍ�(vߕTOl
ؑb8�����ǣ��O�-�ڕ�_9�OGC\�_tB^�o^��_![g�>cvЊvq�7z�gM��J\��Z�AN�=������-.YK�ZV1�G���;w4<��?�9��i��#�bo��	�°g>i��_�-��w2y����t4�@#�'m����H��s�>�E,Y�S�L��K�J��*�c ��D>3T_��***�
��W8�c`2)޳"�@���n��-�Md�������Y1&��̌������g�͖B��;���n��:M�o&�>�sp(�~��@
�����_�z.y�{ Y�X�	�䠲�њ����FY���FՒ;A��#2�J���Mda����5�w7��5�$000�GGR���:��nή�F�?��Qf@�Q;���OU�����{bƱ'�Y��]�|�V���Ό���,��j4	C��?2��*%"$�;s*�a�)�ؗ�G�>��	��e�C\��R�s�=�RI(P�]N�z˽m��_5����D����:�>/�uf?��{BQ�����E-a<�6��>��?�?��u|�9Z����=a_}���}% ��^��>#�f@���%�1�3�rv���QXQ�,$��fe@^�W1{�>5Hcٹ�BT���P!;p�3 �i\�V��"=��P:�3IT#D\\\_**Ї��)Y��D|k_l~[���


Ԑ�����"H]b���e>gp�"P�d3��mF]S�z���Y�U��gE.kNA��+�v����ZV&Α.I�v�(e���BDDMR<e�� �p```�pi��
��o-�o��Ym-/�V" ��:�����X�'�O�J�F����Eb&+����/A&�����**��31)L��CH��w2x�ɩ����v�#��؎ε!�җ%v$�HI,k]h��Ob��� �s��E��S��=R���ԯ7�R����������\�x7�cE_�^E�߾��������y�F��o���
��I0	��6j *�Ϭ��ef#���ׇM[����p�SL�C�2�u�m��>z���#r��c���T�y��29�nb��+H���A��in柞���G�#�*L�`p�LJ�7?���e���UӉ�1Ϟ��R����]c�BY���,	�f㼺`�dm��Ey\ұ����]�gXpQ��E0fX�!�������Mk�8�ƒ|��L8Q�� v�xд�_�?��fQ�3�m���<���LJ�;�|�1��o �~��5���8/v�z���x\������S��O���L翿��������
b*:;A�xd��Ĵ��nU&����!��w����_���4k�M{&��#}��Cs��x'�p��m�Lyfc�=Yȥ�r��.����[��?Gը����6(��n���9H�$g/Z#YZO���Bߙī~.}�� ��h3i^���i b$�7�kW�.��3~~h�n��R�2��z���1�"wH ���{�¾Y��܀�c�CyfbF��&����-��?~��h�n�AؘB:�58�Ywmu56>�7����8���Ň���hw���e�f�)�]�HX@�x��х�T-�V[̨q{c_=5~y����(�?��,�
�I�þ����ܼ�JG�
\��P�S�(z{&�����,;�h��{;−D(U��=���X��(<�ȳ&}f������ܬ�5#��t/�\ssq)<��)N�����tQ�M�zn����w��Ķ�Y޳��6�T��|��4<'ze!�:2�1��`���4{O�X�= ��}��Tk�c�+��?���[��&DO�W�YD�̽�퍸 �/���Ig����`��:�pu�]�����W�U���Q��Ǯ��4��,d� �	砥�9G��4�x�b�H(h��&���$�^(U���F����y�$I�cPkO��S���s���m8�)�C�^*+1 %L��a�!K��EA2�3E�����p��(��2��y"��	Bp+���-�e�EK^Ș3D��cIR�y ��)��1Kԛ�dŷ׼��*��,\��Y��d�49����E	�.��J��0�����\�`  �7]h8�G�+��W;���	�0Z,�4H]�6[��f-�*�2,��ի�/I���ǆI����$D�έ�c�g�,w�^���Akm%�GrE��׊�U6����ճ�v�t������-++�������x���;������{zz8���*;m�1�<P
�a�]@��l��d����%�|Ez��+p����Zy�r}i�H_C��xK�D�(dX?Wt2(�Ea�P�� �=Cɔ6~wM\+��q@��`n��������w�)�A:߁ȇ���t?#`�}����&���]���<�ô�����Z)W7 ��mF�[yO?D�mEE�QD6��)hi�C)��f,]���;�B�%Bw�y?΃
S��Zl�sێ�@�/K����b�P��I�@U�7f�^�>ex;n�Ȕ�!cS��	4�7�B䇺;pm��Fr��d�ٻ<��3؛_!1Ts�ll��̩B�yZ���5��u/O��ڢ6�*��1��GIRbNyM8/��p����\tLAL����5�~�3�H��ԃY�����z���q�t��)�����+��4�������]���䤖F�o¤K\7�0��43錪��K� ?�B �μ��_�1�?h!�^˶�6��
��.&�����F��Y�ʖ/}o� 	��;��������0��!�()�L׻�߁@t��r��)f��&��ֆMq
�ǻ������so�̂�an(#�������	9)��n��Su�����^k�N��$��'��z�j�S�4u�g\���H��	,�0��HMB���GH9d�j�g�,���ת�3/�1�_�mk�wʼ`�C�TGLC;b����� ��{W��ug��C>��6s���x&۷�Z���ON������"/�1��κn9��%;��5��z|�>%d��XHaI)���6��Yj��������15���Q-@\��J�5X1:x�������L�FAii)����f��~��U�(�9�{��8"%N$;��ѢM:ǽ��9%$�
�3P���UR����_!ߝ"h,�s�4<�d����t����~�����%��%�|��_Q�:��D.���	��:.9v_�_Js��
TF�~�ؠv��L�P�"_D�pjV�0��|H,��Cڜ͎��z�������q���� ?�!�������k��KW8p�ox-W�֦7�{;�8d"G΄�2f��|�k_�Q�毬�o�)�$$\�fnE�ԙ��k�YW���)Z1�k�p�����ي9	�|F\��N�u��*K����ܶ��~�؇��7���h`�	W��ӑ����P�yPq�UFA�->�+C<��u'��ۈG��*V���S2&%��ɚ�NZʆ̉�s�*�����Y�U�L3�����L��_�K���l�0�=��/c�}��˘x���@��ڎ�K��{n/���ᯪ���B6H�'A,�����BA��ߔ�o��r���p���p���śY�,5vΨ��㤘8;;9	�{ �G_Yq?0SH~�t�����L���i�l-�Z��[q@��C�Y9:t�~ӽ�4��М�ן|����ʙ�����/0�u¿����I�J����5$N��p��H A,���A��ɓ6�E�����L�hЦ6��H.��h�ėH�T�arq1ryYhwL�,�"n�R�S�M&с��b8Li��QD��Ks��9�q6��SN�uB˂@��'��5�x�F���6�J,�fc��O1���K$Ss"~0mN��,��5�a4�i�&}��ᦦr.�/Ӿa��i@�g,���yBB#�4[Q(�:�CI>��:�S �G�ӡ$]����F�4�P
�5�蛿�ǉ?|��Jq^���W=�Y�8��"LJ��x���l_�5�2ב�3��z�	!+۱rX�fx����"Q�趸9��[�Z�*�P��ͨx��Ge�PX ���,F�?����3�%R��@º��Y�<#�ka�̴��Vx�V7���;���'��������zV.pA�T��[a�&�5y%�P�la?�pF-V-�����(��	Ϙ�d��e� #Bo=<�:��Gj�����W5tXSH�]m���Ts5�J���}�ރNA���#$b0!���?����g�:ʓ�<=���"7#z�`{K3:ԡ�#�=FS��� 2[5�N�4�.w̅S�q� 0��O��'o�k���:��T�/�9@������5b�n�&@�:��9r��^�:����PPۇ+t��
�y�_�@�:-���m�ZA,�;�5=��+�W)LjB��5&3�X^���w�j�:�l��
�Y-ܝ�����4I��9��-x*+I��B�q���DA��O�?%e�^��v'�a$@v/]�;,�ʯ�J�o�(0�ʃ��5�	��T�����@	ǌcw#��hR���H"W�X,�a����[��Is-�ƊȜ2���Qi�Nv�Ci�W8`�L.V�J�a��	Jvɏ��C޶����f�M�qȫ�,tf��=f��F*�E*Ѩ��������'fgC���[�$}}Eb�.^!�.`E���b�3g�����ˤe$���e��4���S���#�_��"�	[D�NGZ�.�d�Q�H�Y�%�)NNN^bW����뙦���@��H׊s ��.��e��]��!]�j�������OF�Rz��i��$���ϭx����J?�VD���Q�=���W��%� �!��!��1��-��())�t��]A&��IW��3�K�:(<�R���Q��_�_�Uv�~� ��d���Qv{��)N,�{��3Ƶ�u�Z�a���'�k�Zr�z�x+�k����?�o{Q�����Pt03BܘR^���y��cJ�i���H��s��� ?�=�oo,	�aM�oZ��K�v@X��(���e�ۊ;����tk렐Z�9x��C&oVH��#�2�Uيc{Ӌd�*�	��o��|ᠣ�z1�Z 3���>��#Fra*^WK�?+���w���� �)�S4p�vZ�۔q�᚞GԒ��Gܿ�����_�P����l�x-���=Q��	���e��Q��B� (��B�K4Ѫ���'�3��-ݳ����r��(i|��,�|f¨����������B!}���&��!��ϴ�.���	h�3�W���d�d�d��d��@Sww%���CI6�`?Ml�	�K��2�ߛ0���Ɋ�Y�X��.T��)/���eP��#<��1��2��!�W �Z�t��÷T�z��%g��bZkE�o$>7��������)_�Ǒ�+�O;�1^�tZ���[�
��N1�9U~
�B�0>�<�7Wd �'n4 l������@�4Ux�l�p>���x�H�������P�%���%|�,�5 ��Wc��+*W��>�����bF�>����}�rcK�׭w9Z0{�����H&y�7�-�V�p��pc��m�x8�jy\ޝ��w�d8��L.�s,Ч�~�@h^��4lϕ�a'LP�ճ�}sF��q�5��"�,��c6YR�z��fnja�r%=(3l��B�n�9JVe�q�)�J���m��C�ۦD���쌏��'Y����^ /���u����f]Q��-�+��1J� A��x���?财���1��d��rI���_� �ʹ\��\c��&��8䌬w�G���~���WQ�r������ ��Y-�2 >·��U�*%?���X���P�a��(�/N���&Z��Ac���Y��PEU�R���Oo��T�µ{w*$+�J~� nv�F��Ψ�+D�`�A�	�G�n�)�UQ�ht~˅9�䀋
�t��I���1K՚`�!�`'� Q$���Ϟ�#����<s�[`c�'�Op�&i�	bø��(��(~�VS�X�O��b"�0�%M�K^��ʴ��S��U�>a^_g[В�/��6��D�- ��x�l93�����PA�9l�+)>��z���`����g����[�k
�~օ��S�Cb_�����7"YPF���kcb�h��0[<P�嬉�n'��8����;�/d�c����b�z�NP��ޅ-)�r	��I0��xi����xX��r�s��>m�����ε�$�DD��"�E-J�����;�Q��D�]�6J�ha�т轎6�#������>����{���k���Ȅ{�g5�SÚK|����y�'�no/�遳&J@��*_�:���1�9�v!$_@�����!�J�d@LQ֋�w���� U�i(��r�lx�M��U��p����)�%d��V>���K� �O�;>8�TC��b��\��$��9�������7xy�c��"Q��d5��s��~�A��-N��LN�d �IR���@�NS�'��������ׅ��l���Y_� �?lB��yw�^�2'*5�(�Ց��-����ng~�`��`�p �T�� D�-�,a��"�Rs̉�IV>h��6����*�����!w�[���bx�a�����}r�{z8I�$����
 Ʒ�Va����o�����ϯ�k�䳉ט.f5��9���, !���A ��!�	Oʇ��ĸ;�x�C�h�z	m�]��5܅�G$�� �=ȁ`K�Gu$^6���S�R�Y�E�Y����Kc�����I�t5���L7"�s/�W4r�?P��3�`�qO�f �;�C�?����e�P qH�>ݤ:%���ѷJ>q-}.}�M�j&��r��[�+�-�y1��Q���O/r����L,�|?���
U�;R����q�Μ={0(i��t`t���ߐS&���&���ۍs�oO~�"�� 
A"̀��w������\^G<K�y!�\6� ���&���>8I�~L 兵"�XU�h3A��<��@U����ZV���H0\6��Fdʛ�Sz���񄫣ף�S��9'2�W�^Ú�r�ԥ��u5K_��Z&,�-��������M?�}���?m�S���Y�<%�9����vRki�g�Yw��|Ի��%'!Clxn��~�m0�A
Plp���%�˰}��D�
��oV�Q��H��ER��Ҵu��
��K����{�
�r���%$�]ox� ��\$C�P���1�,�,�R�q��@#h����O�237D�"k?> n�9�x�PXwT��¥��%�����I����~�[�3�q��6%1p~4�[��":1H�K�cL�|,5D&��T8��^G�*�ǟ߈�l���]~.�b��p d��/��w��E���2�|_e�Ȝ�V\�d�`�����g��'0	��Ck
se�j���7���,ֿ�o'*F��W�P�WHѱ̑�޸殭f��N�.�+���H�>��h�s%F�u�	��_�d��+H��?A��^ה! rZ��,�2�(�~��ǿ�3cus��o�T�Ix{��$��r���^+����p��#����呡�1J:��;�\\�H[�{��ب�z��
�ai���%<K|x����7D�㼚���Yo���#�)��U��:�>�ר�򏁐�zd5DV�#�)s��}3���+b�~Ne�35��)�������v��zg����Y��1]�k�{�)���mB5f~|���&��T���#IL�X�mH��l��OV�8bCD��3;����Gt���<�T}���{���yg{�Ckts�~��P�%o��ǎPV����	�%xG�s��NAI�i�e_R��!��4�)Y,v~<k!,��1��ah�ښ��a��ge��������)� ��d�~T �H[����WĹ�SƯ
 b,k���BDpӕh��.鋵�Zkx�C�ޚ`r!L��m����q��ǶFr��^"D[�⌸2x�%WnH~l������Y��{�\��o�J����G�ZJ��\�gɅ<~������UU�h8+.T����}�H(�� "�$�L�n������r�9��+Sׅ�`��Ef)��׭-������>%do��@�x�Fm�s�������/��vnY}�	G�R��pi�r䘂�s��{��g�����?�7�j@�<l�ueN��\w
�������uV���m��a��k�����D�K���&�i�s:�mp�m�A$�T#h����Џ�7���À/��p�&V(U�2� =F|o< uH!�IQ�����k�W�xs����A����=dD>^�,���`�P)J,�}�I�^Gۈ%��	(~Sɞ��0ᴑQCԝƀ8�p�/�tNǖ�����[Kx�:��9�Β�+���u^Ѫ��El�Lq�A��w��`��<�
�,U�8%T�c�8����ӘG�+����%�jM�L�;���t�6���3�---M�U;�u��EyMO9@��v��i�L���������,U臢c�	yI�1�T�����¼��l� R%|�4�4��һ�	R�,|��ܼ�H48��a�����DȬ��vi&���z!�_*R��~�:��H�5�I���0�aJ�	�rΩ�n����h�����y���u�\�Z�D%0�6د�US*0H:�!���4�fn�Cv�����'<�=�L�r̀6V1��uYh�����X�� ґl�Rm��B)�l���q��<���įN̨�V�����|Gl�黀zp=w�u��n��+[�^UO�uIV�U�qR��o+J��O�P��e��y��c�y�l��τ[�Ʋ a��Cϭ�=��e��z.�����ZN��GN�u�o��Nd�ʋ�Su��U\�����U���� ��^ ��ஆff�<�� ��K�UB�/bw5Oϫ�u�$KA�g	�w�TR��`6a�+}���V9r_���
��S$x�;�����ؼ8���8Ċf���$�)7DH�m������.Y6�񽧱LŖ�{�����Q�zW�Uz���0��I���ҹ����i��n�'�DT��c>GIj֓�W��'@J�k�iĉLjp�(���yo���C~�/��H)qh�bp˲���q����L�	Li��U�n�_a��F@��M$���9�"x��S�|o���iL8/���Oۉ�r&�t�L{�)ӕS�m?a�'̃��-�𰗧�Bh2A;R���k0���:����VN��g�U��B�R�+7l����V8����x�p��lf�h?�o�Xv}��B��M,Տ6h�$Wg�}+W�P�~��yˉ��vPK��G��[�����K��X�����Qp�����g����H�޵�#��a+gF�����X��jݙ�C8���ӒZ%Ͷ��;/���U�j6��9$Y�4،<xv��;S�0}�iW7Z�A�𓄈���?�KZ���7����kң��B6���z ��$S�xE�U!�3��w�8����<»l�	{��5g~���[%�����ؠt�e��G�b��&Y�+�Q	/6q���66�7v^-m��V�ӿp����n�x$��ѕ0�ל*�HT���g>�I`J$E�����un�x\�n�BK����cޮ��PH�����Z�f�v�.���=�UP��'bA�48p;?�I<5�-Nт�ͷ���j��������$kg�?�Yo
�yn�W8�g�l<�#�k�K]
jrn�)�����������bq,X*,D���ZYi���Pz�4(6��]��I
����b.���{Q���E�*��]�����+��{�/4ǡ,��>'+6)�N�S6�y,�}a܎8�v��b������ /{�8�p��$4��w�*�g�i�]�f!u�d=qi��on��wMI垝�"9���$�~vg��[�G�m3�k�#�$H��]�=>O�T�^���8r��j�T�&z�zϫa�cz��:�ƚжݧ0�9�!E�VǢ�"�Pwا�_%�KI�#���X�ٿ����r4��hߑp��5|�3(s�N�����e���[��+��dL�:�3�\�?E�����	,�J�D�Ӡ@�QK�x����WH�^x�6jإj����G�v�����E�b8N�OX�3�(�q��2��D�K_��pvRjE�d�jQ{_T�74�E�k?|�ΒG ��7��ݵ����DG��I���H�S>�+0��R$�D�����d��gg�j�ƊUh�S1��<�z +�&�����D�=�֢0�_������o��U?ܚ�D�S-���L����d�` >���/�Y�abM��p���C��c������x*}#B�~���Ձ'���\�+(t����5��������P�S#���3��(��
j�Z�D�9V������ޑx)s8m�������
�������`�7�Ӣ:�b�۲�[��{#[�i߮,i�iʬ�^_�%Я7�3 ��!��B��UoYU3�*���,�y;�Ǉ���k?��~~����{r����	��w;K�vC�����fp��Ș��E�¥�$X��)h>vb����A��E�l�ES0E�7X��˹�O#�D�����I_zH�I�7�R��MS�y����yv����B��v4-0"IZ�5{���4z��2>DN�ϯ��O�z�f�G�~�=�:>�:�F{�^}|D�sr��w�#W��)n0��Z1�E�}��@L&��4nc^7����y�<�Ȧ{��B� !�(F��H���Z��"�K�9��.7ݽx4Sg��\�`N�ϵ ������ՄƁ~g���C/��WS �X�_+ڶ���%&��ү,t�7��p��%� ��Z
�ri�~�|B*"��rP�Rq��R4j#�1f{w��W��J��~5f]C��k��r.~�3��2��z�Z��?����3�3�m�.��Ȱ���C����,T�o�#y�2��@��Iʺ�,����j�Ӡ�g(*��l�D&/<F���H�e����|(��3�;�{�gY����]���n����{v�T��~��k��հ�!�!��t�(3vA�;�>��H�s�=�q�2��a��Ej%�j�ޞ/ J�����{H�5q�r����;��X����d^�霷?�e�}	T��x펬LtZ+%�i#���0�D+ekN�e!/���EL�n��,^���4H�'�J������F�����M`��yw�Κh)tG4p����(+#*��E��J����E֭*��b"m�Fѹ����h�JzI���	4mԝ����� �>>�t��i�T�&��*��KbS`�r~����v��p�⅟kv�Y$�m��#�m�ݟlm������9{~�����R�����1ϻ�;-�̓�	�ͻ��F�,_�K��_��;�fm_�.�f�|?0���T����(/'�d��|��3� �~/,�k^���	K�����}\`~ZS\�Z�~���K�iu�~�ӏ)�%#}س�` c��@*�0�K۳�5Y��2�Kj��0th������$QV+uUuW�ũ6��)���1�r�}·~�뇤�/z�'�c�	s/~wȔ�*!@6���C��n5���O3���y�8�ծy�ó���X^^nL�
HqV�b�F@��x�jKK�!s	��'�������g�����6q3����O�|�/�d�G�ttt���(���ٍMf�&0ڣj5�j��d��ϹvO�{�i�C����Med,e���©II��Un�=���]2���nԽ�p��l��g�/Y17IF&��IePx�g QW&�;�����'�a� K�>�F/g���@��~<�Ho�?l f���G|+�$66��U�G�Z��
�9�e/�vo�ud�61�_W�<�ݭ]Q�눿PTzz��B�F��IH��P�r�Su�����t��?�F�Ww�t�U0��SB��tl�gW��+�IC���qE˹�LX5@R��A!j��{B�"ڥ{�n!$��%~Y�F!$�~��x���-mp9w��s����8��@;pQB���|S<����G&��e��avE�;�iJ�gĺ`�H��W�۳�r��ץ���I��}���ˏ	�i�� v��`YX�B_�4,���,Vg	7	W'kMp��#`�<|wiip+'ArX`_eD�ش�W�vM)G�+;J0O�}�.�`��|vDr�U6�����(Fmf�ͩi@��#�vK5{��*n܀ԑQB�L�pwo,�E��1G�f,9�[�}���)�M��4oɿ�.��O��s�w�C��K�ل�"��f��$&�s�{��*L�e.:�𘅼��7u���BS����U�Z�8x�4�Bmv�0��;ڀ���#�6�����ￆf/���7� �x�[  �t-o@�cq���U�q�d�8��]���< @u����k��n�$�_ Üs�Û��r�������+攝_���eb�k"�/�MP_.��]#������H匓��S2�����}I[[�{������T���`/��H+0ᵅ���;�S�E&;�J�5��U!�9%A3lh Z����:-&1[�T����[hH�ܜ(��^� ���y3d'ʔY���N��=�	B%n��(��!�Z9��t�m��j�$|)�/�L�7�B��źz����=%W$$����2�@�>�M$�Rd���Y$�rJu�x堖��+#�49��Fj�z��y�l��= X)���^��"���OY��%�SpBm^�o�j�������+�е��\^���E���t��W�8�fu%��=�Ԉ��S�l��l�Ŏu��2�K�%�	<y�|��I���?�q���RVh�Ӻ�+��w��2�dHh��E������\*I���S�ܒ��C�ڞv`K��t�H�H��A�E+�Zos��������S�<[����nW��t��Zp� �z}���}Q,�(ϗ ֩ۄ���(�3R�_�eOn�4�?�TQ愠�_N"x�L�Hu��J9��YH*ć}S�dp�����3�O6� ��`�p�h`p]BjY�P���t�O��xI��I��'����y���]��E�:��VNo7�2�%=qu���.��B������	a(��W�#�̊��@�Q�����(�e9ۡ�yQ��h'�@�\�`ޝ����s&ƚ�@��W7t�!��ק�r�A���]�%�nPJ���S���hK4���1�/��y3X��,�I[����Vcq�mq�Qc�ת���NVv����J�S�~�-��H���T�a�A�a�^��j̜D��Gb�\�+�����%3Ͷ˫�y����RfN�:7��#֤��9'���x���ɣ]������̸�|OiCO�,�y�h7Ck����#s��sr�$K�]~�:�_��~}��� �Rvf���g������i��l����v׹��Z�Oq��+�v޾OW%Ѽ�z���W���wL��a9�Zws�Y��W�����K���f���#Q��#��+o> c�S��)r�ۮN��pb��h&It��$���ؿ"��=:jkBK�K\�[g��z��^�&�mP�K�H�sB�d&v�<��m�v8��t(@���'S�8���L ���:��*���H�Tڒ��+-�9qp�͹�V��$=Z�I�,��|�<���t Q���p�_��J���ěK�6B� �EE�>�lki�#��kfp�V?������ߴ�)��_��u�s|*!�uj p�#���/��B�	�g��)��n�P��ig�3������������R��@'A�FGt,�@T�@Wi�	D�\�E8���hF|���x�������g�s
��F�s��ue�j�.�5ִ֞��܃��&�V����/ �J_��6�)⟬��\}G�?���8k�!���)O�@��[W�RJH����m`E����ޠL�ߊ-��	��uR�ɜ�¢����3��ka�\NB�ݿ9�ɞv[�!�D� �{�R��ǻ>�5Q�.��s���|����!�<��;�_�#��l�9���� x�	��zmd�ڨ�ċ��+|(��c�)�12��"ӗ ���%���uL4.�9@�@�>�=�O��M;�d��V�zz��k��z6��=��"���Sj�O�����Y���c;�	��J�R���OLpМȈ�- �o����5��=xo���cN�2��{��"�ӱ�p�ٚ����|y��7u��w�){S�SHvx�L�<����4I�h��)����U'�ojH�kd�?*�Y}�� �h�i�ƿ�{g�ÅM<���;�=�8� 5�!^��}�a�$L����': �%�&�S����f�u���9��C�9G/r��{H	S��^���쑩+M���Ja�/�^�yr��nOXܫ�4\�H\��ϯ�Yð�)�<���L��O��<�~���!��?�h��^D�zs����N���kt�}�9,O�";�dL��2�#jt�܋�;jXd�a!�|����sCD���M�*A��N�}�|�`���_/�"a�»�e�0����v�Bc��Tc����M$�g������WA2�ą��/�q	��)L]�P�p�J)
�e�y�^�g�^�?����ZY�f�,��i��������܆��zٳe%��������_�� �M�;)O�a��1G<�f��>I"� Eל܂��ã�g��Y�j/�S�wW�u�7�t�H����ιlT�-n8J)�?|]��}T�}/�ѥҸ�Fä��¸a"�0�˶)��9rɹ-����<>�~)�3�K��礑T\S�+�����]��"�(v�P��^#iJ"�$"30GK~2k;�5]&	����*Yu���^F�����d^T���|��H�ۧV��=oO��Q��XI`)�k:��V�G����Y6�.�Pe`�Zd�ZId�ꘅI���U���8�_RR�1"�;N����!��b�nI�{��x�=�L��������0{ִ�ɧ'=�������2V�,���?,]��0����\9�Fam��q�?ZfnP��c��CT�qY�5Zߤ=}�7�q\?n<��A/=+2��x԰^ �������}b�Lf�U���*�Bv�L);�Z�Y�5�ji�p;^�	,��N������(��C"��z9�B%z�mu���,,��\���q�>�3WqU��2�������j~2�YLQO�n�L�̆����"J����J�\6�AB85Mq:σ6Mc�J��+˜w������5��TU��،����!�������m���gfh��[D5��@N�~�1�#�ןD��o���Dw!Bs%d�s,a+�����h��@	��Eœ(���r�R�7�>�T���#��:�A*t��fr�Q�*��ścFUa�͹��)��vm���!f��̥=�ʽ�Yy�
"��\'`��NI";��~�e����v�c�0���#���Пw�~����8��,- /u�$]����؈�&�I)N�1�̪vЭ�U\ Qҗ3�(=�hկ��(d�t	���o�S5�z)�r���R�R"D=[�ۭ˽�^���3�4	I4�MÔ��y����W'���^.hfg��;���s�����k�y;�z�b�/<���'_�
 X$��wL��\d�W�y� ܤ�C�A<�^�Ɵ�s�]U�@�N/��s��5&�D���Q�J�Ә�.ȑ��:{^~������F� DeM��n-�9���r�����o%`����Y��I�9�w�|��5-�$�**�E�4?U��ib-B�����o2��-�e���<8��z�� ���7���d���K���&�Ԃ'c��b�bF�A�jA�\�M���5j�q�1=��K阨F/S��y֎Sh٠Ҫ���xǨ��Ev���f��r#���&"������i�YQD����o��W4����L��,�#�(�־)|���&!yR��9�z��x��n���co��Q��sEc�I����Nc��8N3�������)����j�n���R��8WcE��#\s����b̬}�e�b��v�Nz�.V�91m�� �qֻ�r�����WZ�<?ڲ+.��E�FbC���Q��JC���۫/�V?>+�����z���ʶ�&1���nfNm_֜����-�԰�sLm�M�SL녚�if8�vFUŵ���k�k~{*�b֖���E����� LJ.Nz*0Pf\^&�����t��ɖ�;=�M���Դc�'�8����5���YF��f�~s[���O����;'�7�53fǌD���zy��=I��ζ(��F�e�Ȏ�=��w�E_1��K���l�>`3�c��'?���1�ǯ��(�ְu6��A#��K�o'�f0aP�3�� ���f곁����0mH}h|{S��A��ݒ�[�9/�����P��G�Pr�����+�/O�o���E�{�!D��������q�
�~-M��s]p��c�N��_��9��8�������g�^-��}3��;X��˷[!
�7_nEas����]d_cs�8�-[�Q/׬����i�
�Pފ
~�,�Ҧ��iD4�4C/b�O~��R����L���I�^���e85���|�QCm���k�������,�k��J���]@.Cx6� ��72��Wrɽi���=4�m�������37�r\��4��dlf*4f�i_$�F0��VO��N��pY�m�F��H���e��*�)&�E���ٗ/��o,G�M9�T(|��YR/�5��O.J�eg�Qy��=��`�"�L*��v�[��WW�F��)}�����#��tJ��.�5f���"����	����K^�)�ń�Y�e�E[����a�vJ�4_���~]�h����"�>ן�sJ�X���.�^����s~&�b%�;
6�I c��<������%�nS.u&@�e�z����P���p�H*�45(�'���=��KґU/oU���}+ KʮpF�7�����Y����.rܦ�%�E���gL?#(Z��7�����=�6w����ȝ�\y�3D���7�~)��9z�6�^���S�Y��ձ*0#x��.w���F������Nl6�w��|�����Gis���3K��$���J�W��us�x!��L����F�f��,WGz�J{3�?�������?��6�D�%�� ��v�n��	��d,�X�~5L��Tvz=5��t7�����TE��nm/�x�vc���y��l����5?���:=b�F״��5�X*R�k�9q:\�]j�q�U���5]����T-�&<�r��ާ�!�4.IH 3|Q���\�.���]�]�#��Lc����� '����\ը�3#\�����^�P���&ڭ(A��5�/�I��jz���w{ZI�u��ȉw��I��5j�W�l��^���3 �ȑ3ӈx��:g����G���&����/�وE��D��: �:�R��M�e�FR�_�Q�7��\�����zp�H9��C�ҥ�I(-y��kg��Y3�C$�de���IL���'�C�� Z�_�N��&���XH�s�D��xD��z���a�$;��Y��������ҽ�5���䏻�Q�l��PhZͷ�iu�����Rì϶i �|�NW�T"1>����ƾS��%�#j+�Qkd��U�`�ข��t�۪��('�W����̰Im�ġ�`�U��J-��D>�l��%+��O��8zE��u����E���`l#�>�6W����fTȣ'���ʔ=�N�'Չ�� Sm�sf��]t��b��\a����T�#�2�{��Ib��)D�JZRȚh*�z�a7�BWf�x	��
+�z���r�}�A�gN��)zѺ��f�ڴ�`�FD�?V��[�\�a8\���g(��yS��--�h��26rr�������(��������Ym�ѳ*e�dv��h[��I{ɨ������\	/rŸ�z��u��'^��t���J��4,ٿx��5W�6A�:��&�*�`�[Q��4%��ڿD״{�[MT���"t�,�*�+b���A��jWP�ӕ5�!��>�H�J{�~
S�h�3Y�.F�$5T�57ؿ�gD�˭��F�5���Z�tu̎�=��$���j��E�CL�N���ᘰt��.�F0�f�g�5��>f�c���Z2;��*г�Xu�\��o[�7�q�Q�6c�œ.����K�]��_�]
�;6�Y��,j�ڕ�]���=�@��6z� �v��k�x�����3�o��nV���e�k�w�l�B�N�F(`��Ŕ�j55%̗L��<ཹ#�ͥ��H"���;ﲬ79ӯn#�J��4<g����ɰ�,�z&ŝ�-���U����Tz�&���3�x~ś�����)z�_�HC�5W����OEO�^*�z���X>��*%���Uva!⺿$��2�b )���"l0�e%��̻���7c�F�/���:{y��O��gE��>�|"��6-��L:)=��뻁^Wv�{���%+�o_���{���!5mb��h��l��bK�9��	3|�el�ky�Z��b�$BV2o	�[y��jD�(��ѻME���W?���k������˻ޛQ���D�FŠj�߱��w�/�w�0)��i�gP����=	�tK�iιH[�M$�JP%6�a����|�K�sK�\�A������H��AԬ�V�ط��O� �-?;���R��5b�ܣ�/(����T6�)ϟ�=Ғ'j�*�s��zM-�*\�?�-:�k[�{��j������3>����4X�^q5�7z��:�l���T+��3����d2\��5�B&�jW[|�Kz+\{smez�2��$��X7��KZ(�����/v[���h��l��q-��k����}�E��������`f�`N��A����\�ppWRe+HM"AC�΋e"��@Frv7w����n��f�?E��Md��3�^��^|�n��:��=���=�]�2J\Z�P2���~q ����Y�׽T�sƪD�f�!����HR�D�URۋ3BZM�4�u��c�mJ��������r.�34�)���[R�~���(ql�2 \�jGӬ�85������;kV�Fg�wJ�߷��G�f��:��^YU����i��k��tB��5֨%`ֺ(N�?�.߶v��/���-;��rev=�jp�ތK}<5�×7Q�8(%�um���[1��=�E�1E��O��_β�,~�?�!(��
��O��eS����^V}��l�-Ϥ���Q\�+&���tGj~�xn�g�� o��̟�ǓsGL�ڰ�0m���_t�&�K���,��A�gxw����N��+V�/fVx����Un�ēY��-[tDzv=�{ Y�W��}��Fbɯ-�5��I��<ǧ�"����e�����R����7�?��7�{c�E#��K�$���D�{˷�G>2�6�C�*�ij�p�-�]��Xad�C��c�?$QGY�(s<�����ˈO�'�d���X����q�U�����S|D�����8�mI:cQY��̼�BM��ب��o�g_Ҭ����-}pۛ�+���|p���*37�.�:�Ƈ���$8ު8�B��X��9�>���|�t�#*�s'�m���ճ%�Y�lr�� Ɯ��3{C�O���֩F������6�4hح{\uHW5�=R�i�����m���g%m$��~�R��s���C���~Q���
�4��n�R�G����L�	*_�."N�M-��V�s����p�U�	��;�b�J�xp
�ZUe�j�}f�/wN?��5���#+�:j�rx~�=��YU��_:$Y�)�8��*�£�@X�����1I�*>���<�w[-�jn&N|a�s�I?M�_��Y/�d�j��3SX64u�����!�燜}eM���^�U��qB&���8�x��V�����3,�Դ͉�M	b���%���xGe���^��ON�MiZͭkb�$�q4�\yFs
��N/�du��� �
8��M�L�q8�X�����zH��3���R��z��e7M�Q��3�Zj����׍���Q�@Rb#���~��ٓ��[[�OZE�³��}OϞ���G.D��kZ�<(���"ݐ,f���4 ��b3I��Em��x��2��I�D��U?m��Y<����x�nizp����*��ob6'h�'��^��I�I寊�i��=�qXX�ĠA;�U�e�\6HL�+������--ĥh��gL�^P§�fc$�S�6V!��?���(�<T���OYz	��Ϡ���t ��j,�����	]����y�)�3T���f��dJ�Ta��vH��GQK��Jn]��FL���".��(�;���׃�y��j���n4Fh�]�_Ӳ�����x����Z�ɪ�^�rv�����`:;v�q�||���˲�H�ll�<��Hnï��]7���͚9_٫P_�89���yZc��M��gԡ�l�>����B��:I��݉�'f�7W{��M��bʿ�L�ge4�G`O+߿�q�Q �����r����/o��"_p�"�&���&�4�S�>k�*��ϔ��MC���5�N0	��Y��Ь[����O�3J,�K6�n��;�������5��DT ������=S��d���p�B�Q�c�S�_��G�ElA�|���b'��e���M���'5zΉ	�&M���ZG�IG����,�ɟ����Z�G"�b~���w�)�,XO���5p���X`�%7�R����+'��VY�P��%���cSCַ'Z�8�l�;�g���!�5.�Va���Qm��<Y��<��،>C��}vA��CC{x��*� �e�� l����������Z�ʆ�	fW��(��}jEE�ZT\;GN���ݻl�
��맷� ��G�����,F1��`V��
s3�� ����s&�F��^<W��&S�$M�dw�?y����������oZ�5��n� H<�L�����G-�l�<�zU��N�ȟϝ�}�ܿ
N�h�8��� �#�K(�^�����N��Ls��D#������8���iN4�$n8E#���R���Y��Uř���U_�4�q>��_ZJ��H�r��J��i圭��iD�S͑�5FJ/֩�+%�D�O�d{�{Nώi�9&E�F�E��Rc�xn�
;1cc�	�m�i<,ad?�h@�	��r���S���Q�}��ȟ�;�����X���3/]�RVFƲ�&��^�gŶ�iw&��0ă�G�-��z��Yۭ���\�SqW�{�߄����G��L�j-�l���UL���>���N�%X\��`��;ZyF��ŌV�:�y���q��pW�?�x��u��h��`��Q.�?�����	r�`{D�^vf����*�E�Y�k7��#�!��.kˀp{����ʧL�~m���,$����ZW$�9�h(�>&N��;��6^U%٣�N���%���-�~�u�Y���$�=���� ��"�����`�'�G�C���>���f.
S��N�x��$b�(�޵�ļ��fMڣ}C�=9}:�v,�O�����ƃGO���̠�)�#�ç�f+J*�b��F�"uJԮ_	}��nj�uV#���]%�.E���@�53X�9�Z�xi����n�@�ѱ[���Qc76��9��*�@��*]\�'84�r`�K��Ց]v�~�lA|ư�־˜Ub�
E(ILnN�_s�����Ƣ����Pm��D5h�E��ޮ�V��i���M�Y���jɇ�zi�<X�w���f?����z����vc�anf�^< h6��ϰ|_�V��3�k�r�(Y�ҋ�J W��?���Eg�O���(a��
dH�#_S��
fý�"ECbHՁN�:��AVL��L#�v��p�Xw�t���֚̊b+ܣ=�31�\�����KϮ�M"�|'�h�g����Ivw�0qԩ%��G}(Z�6#�:��-�q��y0�0��O��_���{~�_��F5�6� �m�^��+Z����3\��lO�� ^��g�t�\��j�dİ��b{�N� �QB&Q�ܿ�I��lS�IP��y��	���^G�����k��D�=v]o�-�c��G[L�ݨ�A����Eb�Sv��؜�GE6���½�����y�;;g;� 4�wE�z�Xy-1-�Eu4�~(�Q��`zl�'-�
X���4��`+�)����<�+�H&�i��4�x�����Q���d^���va�Ƣ^���5ܨq��H#O�)��������#�uPb�xH}h��"g�w��H��Ѡx+�)m�� ��y���5$�l���?~y���frdDo���2^Ջ*3D�S�0 �k0����KK�'? {��Ta���"�Ǻ�"��8��ou�h�!X���+P��O@���&�[�}�;{_S\lD�l>:_��
�3>Ϳ�|r��"�8�le�1{j#0I� �4�k���M�����v ��º,�.�9j���նf;5�`���d�l �2��w����K��mYO������/T>�!�"#���Z�����I
���O^?R��;Rq	��z���mr���7[�ۀ%��?��ߺ�0�V�b��9��6�J#��pZv6�G?����C�`�3ZrPAٻ��I��$Z�#M"<w�-��f(]�����C��0!z�n^�Y��gg�Tc�h�#��E'�������Bn#���I���x4^�(��Nڻ�z[�h��^C�Wo�$X
�����T�}Yv���*t]ݽM����_J��.9*����������eVf�2NY �/<���p�}׷j9��3CӐ�N��9�ɻ�,�0����iX���O�F�ڿ����)��>팆�~f_ 	dSn�:ܪd`vXf�x�%�\!�>�B"�0�����A�R����;1�H�Q�k���cTORB�z��̷L��^nv�ަx>��5'�0u�Ā��lBW�,�
����<�m&�:Q�`��M��g��u힧L:5X=v���ƯN���a���lA���x�w@ߞ�9��:��A�"	��r�X�S�Y1ZaU��zq+4��6(��݋������fA�\�3�Y��.�ftl4��MGpQ>��>h��:�ԘV�k_���׾��C���ON��)�hEʚ]�e���e0�!���,-�P��c��+2�c����c섌e��۩��\����s]���]�羟�r��L&`NZa,���6�յ�?��N���b�����8B{�����(�}�����N�E��uog]�Vd�����%��>ĭwBw_�G���އ��UT��h�Wu���M��D�1��Mj�V���Oy��sێ�3���,�^e33�l�IT��I�|�����/<Q�N}\FOr^ttc�&�������w�Un�G%�%M�m���ѧO����+1�O��"�w񽮮�K���a��U-�+�k�����$�Z.�tT���+�ZAs�`���G1��l9KӰ�hc�W����*���>��b{��2Bi�4|��!�]�"�°���f���Õ��Ϗ��j�wP���e}㏞�P���l~���Ş�#NFM��|�zLٙ=p�Y!]��k'K���ɓ;�[��N�1{u��-������ez�ͷ���\�B�ڍw���P�>	:���n&�$�e���ЖRr�=�A� ]��?�8@+��nc�)E �{F�6�z�8�s��G7�jFt���6>�>�ؓL1Kϒ���:�aq$��������u4��e}3g����Hr�sk
H,mV��!�8)Z:���������,G�/�(Nޫ�44�3����A_�>X�o��}�����?��?{��Y��K�����Ԁ/>�rq2�@�X��s��L*�NK�)Ա{�h�^��1A�_�Aίu��+Eߝ��ɨ$�6��}��JJ�	C}�)�lS��NGEv�=٭������Ab�����H��������9Z�W���h�׮�w��S�ڟ ���RJ�5�/s��k���a�~�s�qYD@��E~���&�F���9�ۋ�-qZ��������//o4���<�ZtQ&'u�Äg{�!�lo��&X�)�LC��JR�t�;��Kn�˫���|7\�
.�`��KU����U�6
N��)���S�H<��49�*��e!�L0�_������z̾6|p�;�
S��=��I_�.���?~�]a4Nܸ(��Q�1zS=�WW���C'��"C�eS�c�F��x���m�Ff7�G�=ğ��4	�h��X��<w��w��E���kȋ���E�;��!�u�w�Q� `\�:چ뱇wo?���UY�P:�jZ`BY���O��qv�Ô�<z�#6�hY�
�ש�D�E�{�΅�0�'��ݴ�m���(��d�FT5r��+`ۿFTs�ΘY�w),r��N��tr�e`<v������@��gܯ��q�E[sJn�㈮��v���-�����=K�fcW�R��/8���^�����HE˳LLPӫ��T�F�)���
�i���%�ǈ�~J��s'�${��\�q��g�L��8�3oD��z�Z��:�Շ�o�T��"Ն�!��0�|`�x)KMIO�0��9���T1*�A?���6��hqH���s��۱�=2c��w^�t&6��⡥(�6=p����7,eufDuT5���!�F�(��������<�U�����v���&u�'���]�MC3���m��%u�-kNɌ�P���!(\=[ÅKa�����F�Y�Kg��k�J�	���.ƏE~�^�1��XS�}7�������Q6��v$Tݏ�M�#�R�����9"��G�=��3n3n����$Xd�j���j�P���/��m��Z�lы��Jǿ�|���Cg�l�z؎���?@�Է���m��y�v��\�G�[�G�}!Sz�BI�ЄL�7��#RVIԽ"�7�k�}�Y�E����f�/�?=�Շd�9��a�D�F�|T��������>��Ј�Y�5(�ittޫ�l4X���"������AO,�PVɥ��da�[^D�{,Ƣ���dW ��0��Qswxҧr3��@VYI(�gs�{T��6, ����X�ߐ��ho�	�/$���B�D�?�oįq,
k�Z�?��7��&z�E�1��۸x�*��3�wtG�����;�S�J������x�c�<[ҥ9�	�i#��<�ц�����`V�q�sU G��0�H��֖A����J�:��C�@�5����Y#Ӳ��Z,�p�-��I��;�"m���$v��2<d�7�/�>U��b{��]]ɱ������hլ�%o�����d�;��/1r���Cr��+.�Ʀ�E{��:� �9��Bw{���v��ЃR,��Z|M�6��WN��}������rk:}�z��ڼ��l����Y�������>���d��߳���5�Mj|!�@Q-P�ۡų;��5�<	-h�,K��yM8��0�@}͟� u>}�)�ME��`P���oz�-
k��:`(ix'F�߫�"""�jf��Ij"M2�B$��/��P��3�J]pC!�#���m!Mf��*g�?̍c1�\ c��!����xO�r3�.S�5��I���lRگS��.��N~F,�*��Sȷ�l�*�)��Y�l����	�L����{B��K�y��a[u=�f$�e�d�&FWt_�-�_|�X��8~Su)ㄎ�0l���B	g�����E�.\F����� C΅9������z�b�r-�RD��o��QDΥ�E��) 8E�b�J�&��69��T��~ź����KiCN��%c1G�<�F�$�ʬ_x��+v⣗\>B��z²ө�h|��� �,ƀW����3�%B/z~����]|i#U�1��)6B6`�}/�� 5����%�j�O�11$������yC����o�9�,֣Qo�hZ��@���N-�N�Jg��q� K
��:w��}b"\�9d�R錡�+߈>�R���kg��h@�|�$g�O��8M�K#J�V<��4�o'�#"�2���KFdٵ�S����L��/�ݦ>��������c�$`N��:���`�[lC�kY����Nظ�O�XMN�D��ҫn Ɣ\ܯs��A 3|]X�髎Y��,���K�&������Α9/}�'�ɭ��ʭ�Ԏ���N�`�����_�}��^/I���ƪKm�v�l�3�k�c�!�\��s�.��KЁI3�����A��2��5��vIy�Y�_�E̫�eIy?Ϥ�l�e�:�~`���b�v��Ȧ��ɵq�� �3�Uɭ�?(f��1�;���A�u�.�Mf�����Gr� s낙��smm�-t�Q����=e��S�%c�k�3���{.���������/{��=fLm��+�~1��9�2�Nc*�R�ţ��o�9� $�i,�#�rӢs����e�{��o�i��&}G�:�N;C�8�>8����G����d��c���ܿiM1-#�_I#L�&�UB��� lk���X�,t��d�D��lh	k���y]v�z�<}Ǭڛs�;CkY#\����}��gs�z=g��EM����V0�٥�Z�Kך�����.�g��x��c��^�w�q�[�*6�U]g�S�Ig���	Ȭ;C�D���?~���ml?T��9�gR���ǕX��-vQ��qU^"c4�}::��[��eɇ�D @�^���Xa�g~�
�g�����H�v�ݶ�N))���:?%��u��zdy��-QQ���`?ۻF�HC}R
=��]�����h��<*�D&wմ�U�Im�L��^'�Q!+�l���cQ���W��]�%1H�m�L�8�s�<�v��͜nk.�� ^ ��B+�-k~t*NWx�~����h��v�.�4�/a��9>UG+W��fz��F�#��˼�,�X�D��u>䜍$�o�up.��02ˠ��� ���4*�VW���k�*&M�;�_u�W��K�2j����Z�,�5Z�VKI��:��ԯ�rWCu]2h�pEs�xk�pW��4�-CyX��۴�r��`u����P�'4
Kj��I�b����`��ډ\-��U�YK+5�D�d�?'H�'�:8�.M3Jq�H���Zq�I�8�%�Ȕ��ؗ6�DӦ�W�k�Z��)c��g��Ք�$�\QΌQ|CN�cV��dZ�b�[|��sIJ;���W ���%J誌�3-��Z�Dz_3ZX�U���n4�B� ��U���`M3T�m���@��yǗ�ΰS�������¬�Ii g�30�@���9?���S�!�`}��\#J�Θ�l~U�B)A]/�3[�߿�j��bP�U0�z+���"Û��Us3��W����h9�+4�����)�*q��A�Pz�p�<p ��*$�r("������'�BѷO/�$(=����GA*�10`׸g��7�N7R���[N�V]�Z;�$277'�F	V)K&��<��_%b-���I��<�c�+qD)����~<�4h��Z/z'���/���'����C.���Q�yG�C�r��~��%)���ωP�%3i"P���!ӛ�d�����������#s�܁V�,
j��O�p��rԳ'{�q)<Ô{�rd-۾�(ֱ�y�i��H1�5
4�I�䎶X+�L*>�hue��i!^$�g���_nx�b��%:}�{��M���kO���h�0Pؘx��J4M�4���kO(n��y3�V>����=��L[]�v�j��z��H�U�Y&(�4_x��� �b�c�F�K��`Zb!�݉F&Й�l�e����|�a4��5��ajV�B�Ky]{�$ѹ����g[�Y�������x���Ӗ~�<�L��X���Zm��o�j-<��[�#;3,w�]���<�~: �v����!`,(e~�*p��R\�'��z3�>�RW7f�g+Qˋ��Q�<������6�fD�<���~\ś��%�T27�(���	.�T:A�ɞ�e*k*�Ů��Z3�TPZ����$�5�ݳ]l�gF���9~5=����V3	�ҝ�E�.� �tbR�xP�M�|��_����I��]J��r����A	�����J��Bt��^ނ��B�`j���dmm0}t��w����^A�_����q��~����sx�~w���2��q$�#�?;��� ���o�s�ƥ����H��[�/��Gp�U�x�)���H����r�>�S�4-��Nv���mE���-%�_#���5lX��~�{/������[������s�m��I��{��7�i��]�u� PK   �dXs!��}  {�  /   images/c17cd92d-b315-46a0-b1f2-cfcea726969d.png�g\SY�>�cAQ��� *"�Q�Q�t�ё"�"B��HG�N���'�(�.%DB�HhI !�?fFt�y������0�!᜽�^�Z�j{�]������^�n�����[�%�n���-��ߘ��I��z�73�u�,/����:��n�Ⱥ��Ս|'zJM�~�K���?t_F�a�ŝ6��<�x������ޡKw�Y����֡�i��WOt��O��3uF�.�?Jh;�@>Y��_�#�5?A��ۙ䖥�R�L9ɞ�*�4�?��Y���ﾫ��o��Wm¥nL�n�k�R[�a���u?�qxS��ҝ����RR�T�"�n�����oFio���?�q�٨�S������ׯS?���Ư�[��Е?�)QAcek��h�o&��쏮yAH���;_ߙ��N7!ѹ�/�m�߻�����3�ֈB٘�<��%�j�7f }�KZ
~~,ۣ��ˋ)ybz������N� �e��A'���ˣ��.oH���f���ʞ4xd$�U�<�o�z�1���ڵwS�9a����8z���J�2���y�u�o�Pyz`� ��b��*o�G�D۳��/ep�cҘ�ܮ�%=W
��c��T��,s��;���#��S�'�4��,�)���\�jR�zK%�p+��5�'x���U��u�G�Z#����>���ԇ
^�x�6<H{��v����"�䫇�Ed��U�+'B��"�����3���O�7�65�_��E����1nZ-Z���Uލq�Nm�ě�}�̦�Q9ec\�PsV����퀴^��>l6߿ӦИG3��	�BĘ�����p�����v	��I�Q0غ���6i/Y��&��7��vJ��x\��٭2z}�v��H�?nP�[�#�-�(�'�=z��z&�l6�xh����/�� u.�d��8'��H��/��m�j{���$�E��M��w��A�7��~[���IФO�-w��$�6�^�!<�l~tyu'�i�coB~b��X1��["�c,C��ň1s��x����3�󽿵*�����G,�7]h�4��f��T� m)KA���~&��G�g���U?�����ų[�;m�|�DF��gS�dD��Ŧ<F9E�d��ݢ���J�����홈:y�U�fz4�&���ھ7T��L�1�C�����~�����K���q迪�_�����6��!�H����4+<���F���֢���7��ߪ�)�Ѫ�dSW�.��<��[ ��)�/��;D�[�Yfŏ%}�z���K��:����m��q헊;�����>P�/U�C&<d��]=�!��1wڂR����-�J��Q�r�>d��E6P:�L��^Mu~?�/�|X}�k�'��6ɑ������]��hC_�����o�	�.+ae���v"m[m����5muk���}&�n=bx�c��l�	αck�~R��'��ǇB�G�������1���R�`�_X!8��7�v>̩U�[.�8r=Uz����ȳ�(���Ll
���<�IKj�~L�{vl��|<�k��E"Vcɳߦ������Z�-.���m����k�#S2ڃj� ��ئq��9����6L`۝��/7�͞L��(�0 �R}0�|0�yX<����G��I͕�v�?�Fr�����t�H^�_qLt��{�;]v�q���1"��	N�����=���������1��ú�7;�ffE΀��`�������B�ٻ�1�D�[�kx�:#��� j�/�:/}���PR�c��t� <D`��5�H슛V4_K�������e���0�#mu����Aڼ�	E�H�a�����7������-2ծ�H�?FU�{���
+˹q�ѕ#2���~L���<�S͏����+ �q���?:``�',�:�����{{�Į8!��܏�� �iC���\���©x�//�h_�Twj|�`C����L��OD}^m�z��i+z�z�P���l
���0g���\��Pw#�x�E\> ��E���]qGd�V�=P��+��:�ds�x�䷈1;j`؏�����O/o�����׺Eॶ|t�C��i��ZB E6{�z����πsQ<�C�;��䐘�V��x�����]����g�ͅ�M�iB���=���Pƥ�C��T���B������D�=�=��I~����:���19v� �;��~tL�o��'���B��!Y�k�c�5��WZ�D��f�܇�^^���8�a����YB�b��'�"�?z�s���P!^�IRS��p�t���6�����=g�C��k �`�A���|��%K�����W�����U��*���
�_������>�'��>��"HO�8���}J)��ۗS>���d�]Pv��wl©+���qݓB��zj����:J��$��	��pwQ	�J��S��0B���w���І�-��(.uBſv���"k��=8b��IPZ��s.��m��Z��iyb[b���fޟ2�]#Ž��!�}=D��F���<%D%��Z�xڼ<B���͒�>J똵�����q�ź��e!��ʺ̘�!�o�%��h��9��l]J�������|�"�U�c�\0�D�=�z���&f�a�唖��F#u�eNY@�Mc��~$'z
i| �k�w�Na܁{�1�c���8�r�)>.޽�kcN6���ʡ�wh�_$uL`�����Ylhય��J��X&M
T�,�.�1��־v��}����^�|�B~ν���3|�]KҦ��2�G��n"a�QY��е�G��Ӱ��'D*%�^<KF`}>�]�F^� Ŷ�1��"E��p�K�Ot��A�B֙Z�������a�w����r��\���8��Z����Qd���(_7�/$ת�f�����jQ���D�2ݨ����E-������)Y^Uۙ�B��nٽ�^�Ǌ�pM�H�gG!��5����O�9j������&���·,"�ӕ�j�w��4��z��kGSez����]�X�̠3�I��l��<��W�o��s��!CQSx��Y(������rw��ˬh\E5��Wt��̓��9k0��d _��ײ-Q���xfr.2��/8�� �<����G��?���]�9f��S�-E������6�Z���/���ʶ���h F�(}D&iKpi�g��??Y+������X ����v���s�ٴP��"�ϥ��o?�`/7�l?~�oJM�=b�霤]C��Zu�c��@Wl�B�~d��Ԗ�¿��Kk����F�����h `VХ��gL븖1��:	X{$��6}"���![}��#h��LŎ��#̞�Kk0��?V�=m� ٥�����o^x��I{ǈ̆3TV�����ŏ�Tz �b�iZ)����<��#��\�]sn�/�`K���2�sq�f9��)�+,�c���F^�Q5�=e��!-�[���q2�f�����g}�Pr�)���Lj]H"�л��隶��Yl9�J�����kj��>����Gr�zGg;B?������-�{ײ�3#2S�$h��d�Y[d�<�/+��qԹ��<��Ι��T�O��ħ���ලl�~֕�6KD�}��.����H����Ԭ��w
������e���ǸÛ� ��؉�1���{��pj���{����9���>L���O�8�s�1�)�_% J�R&+�����D�M���þ=��\"+~���Q�r}�Q�v��f�L�e8��:Ǯp�뉟����f��>���c
5N��p�4u%�n(B\�}��g/@:Q�h�`�piu_g�q輡����婬�?*���gG0kx��?�����s{��_�n^�L5t��6�G�N%,ؚ'tr�Ҟ��S=b���@��1��(����F����6(Vc����Y	���F;j��Q�'/T���Dv+yA�v��}^Q�Ӹ\̓�2�)g�\������&�w�����a�1���i�l�ZKA�S�Ez}H��D�,�Hr�W�}O�E2�R�R!W�X:Sm�W^^���N�d|%?�W�S;��*;�Ayt���T�u_eI;�><7P����ɶ�E8��E�iఙ�a��I�D���<~�Į,=�$�p]�=	7�H<�G�5� /^��[Q�u!,�>~�*nљhΜ����{Ո�nz@��s������W�{���GO��H�f.�������G��P�����^j��NA��N)��X�VV4���>U�gf%g���Λ��4t8:s��?�p����c	$�9��6��5t�䰶m&i���^�����i��.��4b��z�P��
���/Hrx��l_�1�\hoEu�t���+5��yh�8ﮖOj䦠�~��ݮM���Ġ�4�8���-���ړV�QPa��L�[�tC'	#K]8�����a9�؟������ج��f�/<X�E��ZbЎ�א)P���1z��9��7"b3��~�?���~��O�)�	3����dØ|RKO顊ThU��kc��=ϊ�e7����8����Ɏ�-�N^V�2Q$�cʕ���w|؇7��*���+��.J�k"<�nDo>�=�Xf�ȟ���g�5�߫�����L��|%���}���D���]���LǓ�P��+�}c�h�ư_l2]O�� �jH�/��y���/u���`r�it,�5�=�`o��
텳x!�[KT�}L`��9�F����f��ڳ������C�/��r��F�#�e��Ļ�w�ڼW�^�'}A~�Qp�=ͩ��U��s��\�����5Qv�����,R�	�2���J�jp���8SLEk ��L��N��k:G����G;��#a;S4�j=Mlw�tﵶ"�MX�=����)�Z�u�a�E��"�`��f��ڵ�EM�#�$�S >p�����)�b�X�-l���^h����q���| �Û��v�&U��(���
�c�h�}��.��`�G�D��d�R��H�l���y��D�����"{�3g!8�YЦYH^��Z��6Jn��>��9��:6��Ά��0"��,�g�bה_om��蔞z({q�U|�\y��n(��P.��m�C�iΦ�Ѿ����$���}�v�{������9��؞T�b�01b��W��N�H�@���B�=Lݩ�����c��I������U�_w'�%7�X ʛ[+|��,SQM&t�/���/��:��>H|�YMҺZz=L�7�fU���
�_�xE�@�<�՗�Hs@�r�)O���/�rq%��*���n�o:�K�����(��W	�J@I��v�:�[*�V��󙈮%�����;��F2����Wo��$Z��B�~�ҵ��NT�h�S��}���#��(��8�dc�T�_�bئ����4A��$�Xs@�Z��/�&�����e��[)0��0��W1��D��[6�:L���s	�ӊNw�;��� ���r�^�%{�Ȃ��]f☷�/��e}�㺯�{�bR��B�J�p�n�;������U��, �ژm��1�a��ܛB��!��UU���e¸�Z�]�����粧��,HV*�$��e�y�6a&?�1�>�?�N�g.�q:�P c�ѕB�p���B�z=�6�6;r��x5"BpB���⏚��>?55�Y���K�i�aL��CK��f�l��b3�|$��D/��g���  p.�U-��.���E��e0u%T�f#�y�����3���)�V���?%�xHۦةL��t �,Qէh��6p����}���i��@�O�01��>fn��r�vCI���lرs�!���t�[7�aJELє�p[��W��u��8[� �Vy�ի�ln�}�����L�^�2����+^��Tăx�R$�r��
/Ȍ�.���� �ɵ�A5NΘ��9�Q�����Z?�ż����+_�7Z�z�=��`'Ϫ�;�Y�%�K_�yV8Z��F���̳�G:؅Ӳ�聈,��G��φ�g�M�����ox\br+�U 9i*r�-�J{�Xt�_�#��F�Ю�e�kN��,�3�{
2?�4�gIp����]~I��&莑�IK �0p�;Bi�kP��=�[E������w�b��^�~��������VS�'�}�) �_�J�t`�"�[1�9rk7�В�P%[MZZR�T��4��yL���<�Fl����k�������va�鈥*��;т�~G~.��D��u�wK�l��R�b��8�a��������\[m |�֛>o���� `!��S�j;�K���i�<�m)��T �����.��g�ʡk
�zx"�`Z��ߗ>Je�+�0�r�H��)Ma�_��2/��#��c$y��^ݟ�zc�n��8��hKó�"�FN�8���o�$�/�, S*]̨H�l'}��GO�]4rh���<�M�����K�,ܥ�=���n9Db%59�4�F���F,s1����Z��#�L�����!f�<`ʷu�����tPcR�Jg���j,����DV���#�{�B'r��0�n+���%��Ⴒp��r8$Ɠ�ĩF\�cE�-����J���ګW�ty;7��3�:f�2I`�N_�]Wz�vH�p�	j$']���>@X�Ufy���3�C���$�B�	��'zjmI3��
}�a<c�q�;�[CܻC��ͣ��]eD���l��&oUR�=������W{�64��T�ڳU���/MЖ/q�rʁ��R2��0|�h@DD�g`�����F[{�����|t���ő�
4?i�b� ���?K�F�ik2�ُV���^�'�ـ�v��[e	Ω�����O������^ L���2�5⍱�^�O�Ea�*7Q��i���v2����H�I����>�!R��a��87��1��$!�gѸ
e�-*]���q"Z	�^�	ā�1kɁ��f�y��8pi��S�aZ����q���|�fRC�k��
��I�˜@NWD�l��Fq- ���af�}g�(�؝��á�U���S gk���J	`ߌ8l�N�����{1p�n���B���e7�h �]�����Ad7=�<V��)���Mpa�}�Y���E@ �	�,�@G��J=�S.�,�~����<��4U�J#a��o��_sF>V�4l�f�^�PW7��"�R���F3Ր�(Ȣ;�sk�ҌS��7`q|g3/���������T���#)�||��}hޓ���*��� �rw"��J|��et@��aM�p	+��U̚���e�gz؏����y�1Σ�&k�+n���WP��l������y�~�VtG\��⤱6�� ��˕���a�{)fzT�_�y�£-�]���6X�r�ܭ9Ie {r�jP@_�@%[�r�?��_½h����%�yE�;o�\��S�|�F�.k$o�qd:�$����~���µ��y>�A�o��(d��(��ئ���6�୼Hc޹[7�I+��rr!�.��ҋ�˱ϸ�S	�m�(���1%u�5�W���q��Z_[Т�Ze��Aw�jir���1g?���9�B5n�l�~�X`��?
er�q�wLME__l�*�7%�b�7��)J��bl������K(�t4���o�����vq�vqX��aa�:Z�)��%�LP��a@�]���	�����hB1jq�K�X?�+#;r�b���t�-�fQ����neP~���%���L�����6O���+�Z���M����4��,H�D�D�LJ��`��V�~u��!��o
vF����*0~3�5P*�]����f�o�x����,�UZ�>=ųO��F���~b꥜^¦GwNΞl�&�8��Cf���x/|�~v�n5�㎿h�`&���'��`�t�ί�i Mej,�^..)Q@YgW�V��]�w�о���ŏ,�!��&��L������,x��� �G��0�`��(�ab���=#��6���J}c�dL\'�2i�u�!��c�L�4���.�"��':cf�u�=��ϕ��o5���Rh�o{5�"��*\���d���?U����#{.�Z�%<�4���S���㚰�~;�L,�c'�U�����Hϊ�DC��T�O���K����U�7�UM��ޠ$J����M䊗AoV:h"��U "��)�C��
�=)�i�봖����,t��o/[`��#{����\V�")�ޡ��{Ǟ��`��������~%9�x߸ޫ�ˢ�l��K폡��MpH�q���Ucԝ��S�`�z�]���k�b���di�My���e�5����+��£	��w�asw��[LP
�K�6�~���F��b
?I��r}n������B6;��J9�bEf�������u�'DVy��ug��"miT��ׁ�zX<�)^֬! �X�
���,xyV��b1���*9�l�\Sm����)7���6{��a��X��E]��Yhy�kZ��f&��
�Vz�3����*# O�뜈��]S�|v�t@#�d�1ɧ�SL��GT��ޕGQ� ^}��p�P�T�tF��UJi*�9�>�W4��GYȵ���ä��߳��-�+���fq�}|;s�Bh0	
+ǰ~�\����5⒕G�{&`M�O�����@V�@� �J8aq�q>"wc�+�>f��������/-8�)�F�Zgv�O��X�BT�0'5t�~ڸY�"�'��d�/
JS�;I��a�z6�C�fW8F���w*��t�r�a�'!U�"��}��� �4�t����X'�~��k!��P���u�ݛ�n��w�~4]����H�<>� ���r�LEl�P�79tF��>���L�!�G�)
�*f�G������k��?x�QtF���T����0Zgp�!���Z�O*gG���)yD�=_�\�(�nϺ�&�'˞�=Q9�W`#�N�z���w���qF�ܡY�R�yٗ�A���Ox��W&����_��Z��@��I�'3e㬔)���N���)�PGƜ5���i|��EU�f�2ӶZ���sVm�O�lFZĹ|]����%D�͙i�XM�wI�D�	
����F�YqV2���3~7���^�����;�y<�F�ZF�k�7�����p�e�Ȃ���������F��0�5���$�}y�>z��k��c�P��%Gl�+�&㛄�e���x��Ҁ/��;�VX07Y?w�S?jfzb��$�*�)���
�|�M+��Q�xg�S�,�c����X����>Kk��nν^����t��1��р��  ߘ6�<��#H]y����^���o�o��f���Ǟ����)��W�F�2\aK����+yJ���>�P�GF�ރ��玲�an.=Y��2�z3�{t�Hj.�\�=� �N�M3ܡ=[ �>�� �B}���3���;�2/�)2}����.ħ�Ə��f>� 61��]���>�|0#�;����F���fB|Z��D
�a����7����͡�����0m�bSZ ���ޱV	S�d����I���&E6�VH�}U`�i4|�V��8۱?�����h)]��.�s�+�����o�/&��K��by�Y�T�>ώ��h�B����ȥ��K~z�ϣ��k��p��6�� �����PAzˮ�0��N*�ȁY�ӣNiG/�]���y��yX����e�Ǝ+	�f(�*{�Ί�;[VQK�:�����N/.*����G����$Q����;�����y�<�Y(�&"9^%d��C��C0'�-:;�f�ڬ�]��;U�E4A5���6����V�)�P�pvwٓ�YC#��p;VU��S������`3NO���~�sFl��F+���N�ڲ��*��E̜g3��6��彌C/%�� �	_���0К�8f;^���,���� �H�]�z�ݮ>�җ�s�=Q��!=�A�WC�brN��D'�9�Q��ֵU�wZzJ�>c��F�B�T?�����0�����2d^r���uV��b���� �1e�k�>���hPL��_өݔ��+�%ͣ_�t�r��dy~c�P��܊���=��WE�x�l�]7��h���>\Q����v�d�x�k�`Ul���l�ә�0�t�Aͅu�v��:L�R�^\"�;O�H<�/��~ܚm��l���o#�~LF��=��6��|��\US���]�f ���ol�埰-Ev��V�6&�3p���� ^�*�I��<i��~�0�Ӆ@�մ4�S���t�tY�FƆ	i�B9j�p�]�}�{�`3:-4�ҥ�w:��FR��jP�.���(�<�J\���
�˴��J4t��gM��>���ԗF6SN��'�s=j|��r�c��V��� y�#�~*�;h�$B���a"+�F�C�9��lE�$�Ai�ǣ��@�"1]�J&=�r���J���ս�������g5`W �&%q����ץd/�ũǹ/%pZ���pI���*C�~��Osď��^n@l/Fte��a*�pl��x��fG�S���	�>%�nZ���E���Ҁ^7\�ǖ�e���=-�~i���4��!R����6I�R/!=M�r�xl�W���#�S6�6��D(���������/f�S�.���1'b-�R��}���ޔ��긖�3��$ ��z�K�JU�K$�Z�Θ��7\ZR,�Ν��C?�^�sc��&ˊ�_ɲn�U�K�G<
�;�
U_]��Dd�hY�/��<����^�~��M+kd9�ն�*��i�ͭ-+�z�E���"��so��S�9^�b{Չ!�܁�p��{����i���Bݵ�X��,��3E�V��������?
)���d��*ٟ��?��p�{���=E�	2��'fL�$j��=�)3�����6q�xWV�������Xj�vW�*"��dig�J�ς�T��fj!��ҏ!�S8�7m�n��jXZl�g���k҈��� �9���x����#�v�Lio�������(iF,��Ѝ�v����}T[�$���E��d�>/�o�DZ{Y7Y��X�R�?ۙnQ�Î�f��x5rT��Q��rw%z�6ܫ�p�Đ͋45b������*�G�em���B�;�r�`:��}��!1 ��R.��o+�&���*ؼ9��N�M}�*®��Cs��9��кw�������{m ���~̠���_�c�rwJ�FW���/�PG�ZQ֡�%�I���8�2��d�c�� �fu��e걙���D��aS���D���M��
�E�u2+����-p(�g��:�Y�^�l��gf�쨀���(��n�8�H�G�g*�����x@x 4����wW&A���R'��!��z�h��2���������&�o�#��nػ��KB�V:$]R#��P�	��j�i��V�N�",�+�e��������D��F���4�Bc*¯o��4��Jj��6SZH�R�bی|�����S�W�A<L��d�L]dH}%�I}��(�YDb��f��	���N�0!	tj���s�j�$ohUe��"�ؓ]�;Ԅ��x�x�9�����h ���Oy��W"ֺ���9�ZeL7�ۼ�%-��o# !%Ȝ�3��xUV}�����v�Z�o��x�9`C��;N.���=+J�|9���O�M�N�&-�8�r����<��2Ճs�x��,�!d������O8ɔ9�<<�,��T��:��?)<����E�T��Ɗ�))Hۯ#���}x^a9grz�C;ߥb��1bN��8ɤ}%���T�V�F._�A[~"ѿ?l��'@�o �j�0�o
SkT$s�uͽ]9�f��X!l�P@ ����Q���J86���rE?b��o��� Ŗ�_�w�T_��*�I�Rcz�_���QK�B,�:��x�A�"MqG�X��6Դ�=�(�X lRV��2����dj�y��jf1�خׂE=8b��8D|{o��/6.`
�{֪��f/U��˳tӷS���2Y�r ������pr3��D':���*C����8����)�K�0�P�\��K��Qoy��,Bw�t��b��sNf���j�:��֥��,��$�2n!]`*lTҘ�o���}k��"��D�a������FK�
_Zn7�LQ�*x6tϱ�-,�=����1uP�3{�e:��P��|��^�@���J�5�ls����ώ�,�Zz��bT�1AlfR�x�����E5�ƹ�90Ѯ�EY�-;d�k��B�sPES)-.e�P��a,jolH�3��P�3�~�+u��1�['��oR}�D�N�z<-��#Ւ��h�P�7���"�z���J9m�R}8�Xn�/ h�����wo�ݫ�eZ���W`@��[E6���0B��C׌b��PQfV�Ѡ\�%X���Mq���:�M��,�[~�jOX�w����G������t@��:W��>���Z#�U�é�H���ec��lnp,u�S��M�q�'���a`Ϲ��=��o3ǂ�i;&z�Ý���V������d<a���5�S��"KA4��`M����D<H3e%̷��G-�oؒ]B�&Y?��:(�'�fP�T�G���.�����}1�&���rX�ٖ;� �o �*�� �)Z� �]�nsɧP��젏K=���7��ӿ�
��o���D
z�.{��s��+O^�כ����x���ȿ����ڱ��A�ojQ�WN#��Y�6Ü�+օ�s��
��,����`s.E���^E�"�0�(� ��V� [%x͕�Y{"'��9������<����r ��dt�c���0��g��[v�؀Yj,jZiI�ò2B�I�����9C��n+�S�d%��9YA'c��u8���ﺒL���WU���7����߸D@����0��XHP���:�7P~s=�G�OI10�Rj$�
����T٩p�M�w��ʙ\8�aւ�[�;���Z`KU��E���H�_��P�O(s�#���pD���J�ũ��k41�欸�:��i��Z���� ��,|�j��A��)H��&��"��`E(�]�����;M���B}E8j�cWY��������4�؃o��-`6�5�M���,�^*����㶈,2]����f��:�ٮ����,�^�~��/�H!.`���o��k�U���)���E�,����z�#�{/öW�(i)��BO7g�3����#&��3NKA��Z]U�w]5��\��X���q����*9\�OE�i����Lf�<���-�!�x�V8��L��^p�;��Zg�!���ٚ���\xs����aOǡ%��3��D�D<��mp��F=;WM�6�v.������5<2���s��V��傥�
K��v�D�`r����2g����:Ǘ�c�
�&G8�\D���}U��*#�S����{7�����v��0ѕ��Fa��P�,T�ܫai�{�̨Upu̎�we@b����C%f�7��b�P�����h���G�(�J#`NR���d���[�Ĭ�eJ���'�������o�bݗ�w�.kq�@�1_��S��uM�M��3�
8��O} {5��{�J!���xg�b!��1��NK3�X^ˢ�o�˳sǭ�I)������Ơ�N�����@<��;�Q]�n�_xa����І2���W>��E�M+��r� +��3�v0��S�
r�K�E�pF#Nry�^-���i�q�=%�����!����v�7��Χ�<6�$��2 v�u��@/��SXs\v��8T�W}�m��3�+hܯ�{�?���\�89B6L�A�8W`Ҽ�*�s��MfT�^��FMÆhVý����D�"0&���vf�=�tL���l��v;�ѓ�{`��ǁ��u�~��	�v���e(z������N�!a(�"8X�Öy��el�'�F+^��z�Y��Y/�Wj�M�b�NA�8����|sY�d�Bɱ��e{�`퐵i]챏x���]ͪ^�z��k��������d�{.2kQ�����M�@ӟJ��PkkCcR�5�y��(I� Ν�Y���8.�C1)�}ei}����I��'�nuK�{k��.������/r)����,;*5 ��Y�ݍf��*^k����
/���_
��m\�q0R��aX�ߋ���*�e��g<�B���S.a6�&G�Խ�Ɉ��bV�5�����4/�L�=�B�Q+�.�(�h+S���s�=�SP�:�CȨ�|X�Q�� ��<ml����~_�1�����k��$�1a���rlI�_���+'��l���/����ˣ2�8�˜�Ղ���wpox� d{A���+C7Z��U,AN.��,���\i�]$��M������7�/�f1&��Μ&3�W�|�zCL��w|�{w��3�e=.�VIj��X�hv�p�����3�).����WXs{n�\i:��av�JAM�Dk�j' 葡���`���J��<�<<=m�U�w�N��zL���H{BI�K�}n��˴��L'=o)��/�,����C&_�VŘ~����F	�mS�I<z���+��D����[L�iby|��,�D( �w��������L��h�n�SN����j�.�R�T�[C�b��^��4��mĿ|/8���\��ޘ�x�З�z��:z$1 VJ�����ni&[,@u�>�����/����?J){>�9�e�ҺE���m��a�ki6����D���j.wf����"Ku�����XU؁�t�o�f���kJj�>�Ք���K����g;���3�9��ù�{�@�f�,��b;�ٺL}�/Oda�sG��)����I���i���Qt��Ia�̓#�5ɽ�&�l����$�e}�V��?* �B)��etfGA�^p8�^i1��,���N���7ݦRs1�)3{[��[��F�#�����uAF�@���#8'K��Vae�}K.�0�e7�\��n*�2��8��U���2Ig+=�&�\:��ɉ2���8��]F8��Yc�~�ҥ���φ}v+]��ڨ���5������ ܋���?[���o�����n.�#.o1���%[kj��.L�$}ȼ���-�r,An�@]�mX^�Z��	���-��3u��
)=�cGe��
u�N���f�;�п�4s�vu��z���}ZB�i�b��/�<��p�Iv����qh�P���u���O�D�喝۶���g�G-v���h8���I�n�fE����V�`��JC�h�P��8j�N��^ɼS��f��ř���z�%'�������C��� #d�"5"��+k�+���p��1K��S�$�m��Hiv��q �v�]�������Ķa���-I	N_�fk��h�E&�KL�ǹ$[9�ρ9_�dg���I�~�c��X�����Br�\��ѥ}t�����~u��:�\��3Fd���~�U5�#c]�������rx���s/�p�P;`�35Q����e����{�&���*o;�a
=��OyvL��Q�n���{�^�fWj5�_��Y�u�;b���������ъ��9j�Zg�*5�[vd�K�j���7�֚��`@0�#G�\�^�^�����m����ۓ�2qz�����<1�L�W�D����[h>v�Uj�7��Kv7LA*K!�0;_W��Xt8��=��:gzQt�;<�0Oխ��,���L��	���A�~cӨs�GE�%��3���Fe�l�(��������ǲl��/EV�xh�u�{�zb�yT$+M�����Ѫ�N��Pn�)��$sƓ��O�vd�
N���4��D��j�F �&�(PW�5�/�(h�tb�Ӫ���d��8:ണ�@����i�F5{��L{�@"P��N	�ꀡ��Q���9N��H���m�s��$ D�z�H�n�GP%BX�&�d��1����!q��8��<�����\c��
l{� 0�W�{��;L=0�m�Z� +��	�#�${]d��L��.ʏ7�њ�~/e�O�R�]��̞��5\���wɖ���r�y���.�e�雓�� %dpU��a>3�k"�	`y�e��p��3�Rr��#�-oD�<>0��-���?�.��#y<��X�ݾe��J��`+�⯃y���W���G�L��-!3q%ں����z��bU��X�,��[��Z���:@�JlM/���c�j�8e�WS,���vik?�&V�Ŧcf��x�C-���"�9$q%s�6����z�H��IVK�v�p����E`ڛ3S����'�'@�+sWW���ڳ���)  2އۃ��S�57|x:}/�0㱽�w���9;%P.�W�{�����Yb�>{%�@�Y�z-�r"4���1R�؁2C1Ziy֛W��P��_y�K�5W0�\���5�����E�0R��G�S~���u���{�Ym�D�~��,Mz]Vĥ��U�RZ
�\"�7`.�j1�: �\��3�>���e_RUś`��؏[J#�wS������·�$��PV�)�I�<�@��d ����������%�Ly��>�5'�rc��z5��w�����������a��`Y����+������2摠B�#=�ZңN��G���
n�[�p�pLl�"3���GҪ�\�=�z{�*A2ذ�d�/���p��^�r8��(���``C Zm/�f��߻e�ջ^W!���~���\�����Ϳ�F��۵�y�}~k��7 �<��������n�^^��_�F�g"�"([���o������#:n�<9H�y�m5G��C[�~�\��u���v���i�Xj��'u~�O;���^��>㿇���*��e�$���,�z3�yZ�Z�����TXE	����U�M��'m��Ts�~"�ȕ��ϐu=P��㾓��2��h5n�)���u!%,�9���U%Ĕ"��ZqkX�;��*ؿ�p�)ͣ��N�D:2� l������T]�	����,��~aևP��j��6�Yp�d�ٹ?6�ǵ��\4.8*��M�7�������1�'[v�fEv+�J�]%�,8������7zy�6��#2Z��y<A.�y��������J�ϭ�����A�rW����H�恵r�|/*��u��OJ��ۻ����"�Vf��	��7�k_���i�ʛ� �ڸ1�T��h~��[������!_�<K����$�lڑg���f���.�|�#��R�O��w��v�^և�Y�T��ʍ�je�2��xB��	�-n{�������W�/� +�J�s%��5�}�Ӳ$ul�}8��Į�Q�{y5 ��&��|�l�6h/�"7{�ȈY�*��d.| \�,fHZ���Z�k�e�8�����}�F%Ky{����ݰW;���5˧�Oy��ɳΖU.����~o���*�l��E9�xyKV�ʾ՛������Ym�����p�B}8�I��E��έ2y�]!����@�������	"ĝ�I���Cg��E=[��iqa҂��uvE!����r��Q�4m����i�y�0E���(��^��&h��}C������ۮ8|�B��7y�:6޷������8�o�g^���k����H�7^X=�U������Ce�����u���{��̹e����\�-z����Ko?��{hԋ���7%����BW�-i"�6���u�����{�M�%;��C�8���NgD�N��3���]��vĹ���w1�a<��!!���j؇'�0�:"5�iF�����^C�s��j-q-�Zf�fP#��6�b�<��D6���=ev�I��Z�d�����d7+��C�m~���y<�{�\�}r:D˩,1EQ�2��Ӣ$�)	Y� ��e��)[����M+�-��ӡ�`��6	31�`0��\�"u�ݿ������q�?]�1���~?����,s��BXq��}a�7�W �U۩�rŪ=�V��8޵����8>����wy^�j�w�u�u��Ā��?��Q8�7�7�9�o�3�<ʉ4��!���4��K��>@³l
JkL��nj������K���G��5�J]i,��t�i���b;`�h����Qkq�פp�Z�	oK6�̈P��>+�{�ԩ�?81�XM\�$Oǧ���p�r���� ��$|Md�����_U~F�Gm-N�8t%Z����e㡟�1�x�^��/����nY��:����/~G"b�L<)��O�e�]�<= �2�)#m�F����X��]������oN��g��\oG���w��6����-���6̾ن!��G����V����&���Y��QF��w��	[��a�ؠ�W@��7��E��܁=o�*\9�$��F�_�8~s��%)��/-1�M���sY��=�����~�1� _����K���w�]��Nߥ�вu@ٜ#���]�	軔����\�F�P��B�s3q���|-����о_���� ��^�Cl�lї˅���|��^�\�u�Xq�=Q�M�D}�K�W ��V���K_A߅�%�lUЗ8ޞoկ�c����
U���k�+�o�Wʨ�;��)-,����Wo#կ�F�u��w���~�']�.O�:��b/؃�G5?������b4ӛ�eH���qGoWN��D)׬�ެl�V9[ן�e�Gy��/��hL�)�O��X�>ew]��������k��dII+}�A�ZpMJ������<1��>�q2��-�k<�	-|�w~0>>y��ҡk��5z�M���E�1vQ�f&�u�1�veD�> q?M���27��0���2_�z��UȡI�#��]���m*]v.h��@cl��WZ�4$�� �挴*���XVը~��w/y�{�?��>5�^�{Gb�Tm�����@/ѡ���h�����=��;<_�!Pnr�.����L����C���Fn����-�Ĵ�cy���w�:{еIs�E����![2B�$jNP�t���7h�O�?��"Ϧj|�}���z+���z�Nv���Aw2�G�r䘩8
�t2�rGSu�%��z�^�q���H�fq($%gt싍�]�o����Iy0/ډ'8�M�\�3�.�N�z}��јc��{�IiY����m���UZ;�d�Z�k��H�}�I�9���r����3��NF�2�C������]�a5U�!���� �n�Ӻ/��ເ�z�)ǻ%b��V�E��!��Ul����Wz�4���9��mNۀ����づ/�+�}s�4;�n$�Χ-��ؑ�J���ʡr,��o��ZN��=��n��s��_O�]�L;���Y��g�΅�$�,��M��zx�n��MjD���XSVRI�m�x�*Q��t�,����s�=;�c��sKzx���c�Oy���9ͱw+k�ʷ�Iq����o�>��G$8�vw[�S�dj���i�����\G߅׸F��c-V��a���ĔD��,��ͱ��w�Nj{�:�y�z*��j����y��o�N�ℭ@�c+�{��$���8S<bSMO�|Hݙi��}WAʢ�oB���:���]4�����D����~X��7��.��;)���;34�T{7���ɇ�?�����W���(�)�N5=#�2��1ʟ1����w��5�I�9�n[Ny|�]��X� !t6�!��JbYM�*B��%��n�}���ܽ/�d�I�S�m��U�8~�H��S�P��F��e�X0�잓����OZF��dOPl$�xݣ1^��+?�z1Wu����6H�Ϊe�ױ�.,*Z��K�v�|4���L�$I%Y�imj�\�!�>��[9��1�|�dIѡf�dʃ���a0)m���08�V�>�33��S3�ĕE<�5U��&,"�;�vX{DP�������InR�g��K�ٿW1���/�(��FF�d�ʚE��CO�e�_3#p*��tt2s����.!R+l��b�UP�_D}^��T�	�i�fk��Tg�Y~�|W)=\� >�%�o��~n��<��I��������B���%O���+��d�N2-��{Y�d
B��M�e���]���h�EUX8�2�$��7�W��+���w0�1je�W�{�#ۃ��[4�Fy��*�`ř��H%]�u��A�����^Ad�6N���^
Ew'U��f�:��$�h�E�z�!�Yb�ES�j�`N
��B<x�{8v�rC��j[���33=]ባ\��)�QC��v�/HR�T��Jm�ma�W��`�=����Blx�]�g�J�Cb���V`��-�D��xo�J�	93�[(��R%0�Wx��
5��2�E�'Do1�K���?��5 �ٙpy�u2��y��$3����v�A��7���B���V'� �> n�=�Zjb<�?ڗ{�/�>_cWAq�M?���:S׶9��t������"�S�D�N_��~R�,X�|fft�,	�/�݁�2)�|daoI�ߑ�1�� 5kx}�A��!�l�K�#�� �U��N�A������$�#s����?�z���m�yn�� �\���	���Ī��r:X+�/��"�j&F����y�ow�U�g�G?
G�Oa��8PKt���	ƙ�����^=�u���|�v%��n��mP��}���h�c�����.��v[;��#��>�=��*Q(g5�3j,J����ىK������n���s�2_~�a8a5�ϡ�o����Puy�̫���d�ۏ��T�-ܹ��G-�ǵ:��"K��]o�&�/8E��T��O�WW
��"�C��_���x�Z�%�,!�!޲�Qn�i���=��>fR>C�,�� ��P���(��ns��u��2�q�� <Yo��PTtl�`��q�E���	lgݲٔ��  {B��R.q�GF�E�������qLZ�J�ڡ�3�k��۱q��0�f�E�@�#����BH#NG"���E��:���")��	�ai"�N�.��T���� � ��G ��VY�7�Ќ�V"M�	1�ޟ�_�|�U�{v��P,=-ݖ�+[�0~���I��0v�N�+�_�>�I��+����Bܞ�ۤ���K�Լ�m���~���D��z�3d��&$��HplI�Y}3Ϯ�N�6�`^hH�,h��)s5�7�x�Ğ�=�f������^C"�o=�l�;��Q��:��s�" ��o.ȨQ�.�%���یh1R�n�Ffxn~,j����Mdz
����J��4e
P۠�,��7yi�^�ɑv{��iy&��n�"��{?9�&������㋗��:��c�.���ne-x�D�"�B�Ǻ�s�UB�P�r��A%�ᡃF�6��d��	����;�^�S{�����M��r^���53i���L�s�RH[����O�ׄ�O�q����2hĽ��MVE�ȣ҆v��+�/����~�k1���"8)�H����1K$~~���?���!�Zm�u`��_w���"�,�M87�5���a E�
�7��6Jp�`�g���|?Q:^��aE����r���C��i���0�*�3Ŭ�e��z0fv�a *��\-m76ڧM�:�)?���\쏁�4�Zv_��Gw��9w�ֆ@������w\ߴ7�ĝ`qձ�U���� �i��?��7��� ��%=�>�q�Ք��t��X�rX��&|��g������>/^�jcʮ{*9���Gv&�O��R}@Z�{�]�m�E�Z�=�X�y}jql�J��R�@���!�f	e��U�O}�����:�%��O�h� d��r3NŶL���̟Q� r4�^�:�uO��9hu,E�hK
���!����s�%`I���� �]I��f.�|���d\p����:[�o�s��Zo/��=.��Xձ� ��t��7�%{��N�S�)��]����$z�٥$cH�@Ћ�P��`���A��Sg�]��.�Ҙ�R2�RD��3S��Yn}ei��肟�C�9K�Jٳ��̫c%��a�{��n��ؐ�ϟ��c� ��7�oH�>��{�vq�-�_�����B�sQԎ
Y����n۹�!��k<�]2k�|ui����kqRچ��)�k�o�Eb8���4]��Ǭ	R�/�
4r�5�ه8��LT�AB����A��2�A��&�����(��G�)s������_�f�����L���͸��=P���ex�o���@hh�qv︺���mV�se딹@��t��b�v�x�u��1����I ����\�U �T!2vJ	� �b��$*�OޝPIC)��#�Y�FT2�$٣1����He��v��}���1~|�����n�#�D�Ő��E���#�۰
�u����C�v���j�.�{����g�@)��!*�[�|�kK���i�ӌO��'x(�L��N� 0����vnʒ��|��X���,�Wɜ��Z�L�Sk�	���s\���}�(��*R���iC	���s�oT�궪-s#YN�K�h�ެ���na��p�{�,��v%̾2����!�ç���ચ5�K�!j��C��-�Ý֮����C��l�VN�zTO��PE�^��Hʲ��U�a�+��v
(iB%"��?�FC�!�;�-��k��a�;�FSuf�#7��EG/_���A����Q'x���s`NU�L1��`�LZ�y�^V�w_���t���o�fT�
�m�Hgi��z �K�tJN��Fyfp�7
��%��v����`������Xu��]�܋�rz�(b�[�}JY�AZ��^� �z�����,�o�di�����ODl,�?f:�CTO��!0�� >f�u�/�A�̈�Ӡ�a?6���Ҿ����hE��	)�fͿ��[z2q�-��Ƥb1L-�hN��[�xh�E��J;� �y�mF�QU���..�/C��,�{�w����-o�|�"�8�
�hۚ��  ����AϵM�}�|��z.�t�2�sd.�!L����Y^X�$�Fo&*6l��]o����7������x�Oߕ��o�.���)"�'VR}/h8��)���Z������I��<�[��e��T`���c����?˞Q��7�i�o�M��p!8VM��/0�~j����R��QA�* h@GH�9�g���ʢ�W���^*��A���#�ۛ٠�[B��z����Yڇ�(��o�g �3�6.q}�is{�����TH{�v�A��B.e_�X[��F�u�v$WQ�-I��M��c���e���ԧ$�4�����l�RF	�:��?6��Z]kF}�<�lW��̵��NX�U���ow�B4��g�23gj%C���6��]�!��'�x�l�$�l�ոv�▶���W�~;�k�`gf��٩��A�A�������R�É�)3���R[Qs����}CȨ�b��v�3�Π����:3V�j��]�Av4*�f��1�\0�_`쒓7�~������$'!j�)���z�>�&O�đ���b�Z¹/t�Rs��>9��]�<���e]���o��
�h��<a����U1}��I�m��x��������ǃ�2����o��d���m��E��ֻ���s0
_C�J*�����^+Ց�uy����ټ�cW�e�M�kj�Kk���Hk�2�L�+��w���B6�z��(��>G~)`�~��t�z���UO�.�aH��_��P&_zO��:�|����:�$��6ysH �[R�Rv`D��W��G��_�����>1��Nk��?�Mi��DT�m�C���-y���3k���6l]"=���!qV[�KR/-��)��Y�)WZ7�ϩk�"�x�A��ȡ?�p3��̠E'F5PX���mz�~�4��O��AD{���_� �mʐ����:���a��E^����L��i�}�����v�9OI-nH�׋�k��W+�܁��f�=%���e��=%�qB����V���DK�F�@������)��ݬ���M�5܀��M��v�̃v�v����L��=�n`8��t���0�-:������h���ȵc}9�bM��L�+��O�TjUpő��,�}�$�/AU���4��B6����>H�c��\���W4�W�>��z�~�^�q8��n�?-�3eqs�߉S�#�!O|7<��>�T%h4ι���zCY�#��k��O;F��>>�-I����?�e�|�^� �;��������/�{['zD9,<�s
�}�Tr�ʡ4�Xo����b�$� �Cn+��'C5�������ќz���4v�F�k��J����Ʀ��0��z�t҄k��d����-P�~�G�c���,̇�¹��)�HA� ���a�7��m^j�
6�Lǳ,*���=r�b�C��	HVc\M!Gbf7¢" ��{����[Y�� }ZB����D=�훠)����(�d���x#3�5A�*�ˀ�N�Y�jrўO��q����%[bȁQV�o2��RU�ӂbTĭZ��:կRꛘ�Z=ɛ�ό)�Uu۷p?��Tig[ �aiW7o����n�d�P�p�If�Y�6x�}�
��3��A��}2�^-�?]2�6Li���}����SL:��-c^׾�9~S��gNr�&���I}�l��ô�)��(���踵�6Z�4�H��.j�nMt՝f9��J���$w2�h������<�������;$���fٴӓ"����f=?�hG�9j�.�%sWvׂYz>���	��l[�U����0��X9���~�EC$��� j�Hku���}}1��S��۬Z��d%�E^]���Jgңz���j�f�1,�=�b���dĔuoj�MN9��L�I|���	��WC�G�ҖeL�R�t;:P�ϱ�;�PX�d�j�����3�ֲ�{5�h�7GQ��,sm�g���ݷ�mB�}�4�l �Ͷ�<�Pu�� �]M��x���|i�D-����.�C��bs�����+SB�}!G(�W�$<�������h���`�3��U��~�u�a�����6��e{t�"��ꨊ�M<|��{~�??�'=|\��VY��P�(z� a��q<0^(�"�~sA�I��p��L}����?����,�H2v�2H��]��z�u�����L��OAf��H{w�,{\��E�����E�B���ق�\�	�q3�a6-�M�o=<��!����p�	���^�<�z��@����1��hdy'�1+�ar�X�	u�zO���̬���j��!���a���s��:�V��i{һ�PR�R;MD��	��M��L��:K�M�[�&(���8�f��}����,���a;��x_;��_�&&C+�'H{�4�j�N��,FZ2Yyjf���/��p�dI�u�����^��]H*`�x��:�Ȗ��_b�e{^+>����F��O�n���ݤ�������"H7������c��s�Mhi��e}��b���RCD<�0kyo��a��PD�����s���g�}� ������ْ�b��~ ��|�I��p�8�KZ_��ۡt C�i_'�G�P!�A����>p[,24�z*u�$��ޓ�꫟��ڹ�c�]HY��%_�T�6�e���/da����qܑ�V�e�i�;�:Y<�5���΂� ���-`�=�������M�gi�����qx�5���W��Y�ϔz�;?<����㲎8]�!$�_��af+8a�T�%��1�A����=���
b4����~�<�q��Enz@���H�&^I�s!�z�^)��ؠ���,.4p���f�[G��X`q��~�@|۩q��jkykv"O�\)��{�u�Ȯ��|r��rz��@z��i�G�&��-���;)<��p�{���UZ��IFQa����\��忌1�a�y)��7� �=���\�˶�d��Ƨ���]- �?x�}ȹӻ\oHX\���+��\Wt���%?�1����2�%a����͖l5y���b��ׅ6�X6k�%5���ʺh�nY��Y���8/�lr9¨я�8���o�3�P�� �sY���fI��8	�	+N�}��
���?�v���`o��Dk)� ,�ik6��?˸����
�ٕ03��lo�)/��B��ĭL�hO�|���)��Qk4?�Z��=I��Z�����Vʒ�� w��j���~zCƉ��R��lX���%J���ؒ�5>�ަ���|�I��z�؛�2P������sa�C������o=.��mы�� �O���&�鄾��=<���o���� (w�.V'��\:9յ�2"�l�	&�\�.8�7��1��%���$������q��΄��}?�	�ϿmmU8\s�xgVٟ�5���':-�Z=���})OA؁��DvK�6�=w�����J=H�PL�T�3���Щ�SOw�,!�9�%Im����]��[�q՞7�2�Q�0�k�xS�t��)z�)�v�bKHR�"0���7��[9E��#�v,թ�?r�P;h��bz��F�hߜmS�4��¦��ܺoRWp�_���г.G {mP���u��6��J�-����z����1���%fF��+wZ���c�]}�v�Tz�M���R�����b:�*B�m]�s��D:~5���kw	�mփ�ɑ���"�5' �8�*�#� ���ayB��>�&�>�47Y��y�n|��9�,
��*���!)z��2�4FrjX6_M0���C�#�`��d�Ӎ��<��e0��#?�:��.�?,(�X��N^�t�QhYM\*���p�x$Yl�c>�u�4ְ�z
(T쿨5�c	=��W�2̔��x;�����!{SYo�Gfщ�[��P6���|�rU�i�N��z�6�����h��I�]�%&m��������y�P��Y����0�Z Kc����|x�_"�VU��R��f�|��������}\Q�O�\�qY���L�1�v�
m>�)	��h�2�JٰJ��Lu����!�M][L��.��t�LhU8��=İz��ͫ �e;I �l�ԶX°F f�����l��Az�6��8u���A�0ZF��u�Ww,�����Q�$l��~5�_��rPQ;�Xq�x�,�1��%��~F�C�0���!,�Z������ʑL֮��n�P�m�m�̩�k� dPܗ]�ko��Ӂ� �Q Z�j'���UDs��ŧ@�>.��Iv �+��lMy:�����4
�Φ���D���}�ч��+�5�*B^�+^5�HDy�rF�陋�/���Vh�.>=F�W��Z�ُ9�g��]w0WM;�i�M���_`��F�S/@<&/���$�`��vk�.�{�Xh�߾%�L����\�Th�آ��xu(jK�Ȳ����r������R�����I����Ч]�����h5������~�� 	ht��װ[��$r@�XES���b�y#�QmП;Me���#t���Y�g�b��8!	�[��M-S5֮�n.I�P^W;�<46������Z�gJ��G��̓U�dwS��RROW�컺R`
+N+�i�%A57�t�k��"��ϸ� �������xu�^���eC��n, �1I����י�Hrq��2/J�A�W�����@�y�WѩQ�{}(�o;/���;Bˑ�٬ѳ�?,�u��g!8~}�7I� x��s@w��W�%�����܊��.dU�Y@��T�ߦ/��ި�)�v(�jl%�+�
A+-��~Z� no��Q�vq�i�v(4}�d�㫯�ұ��xX�b/�FA��}wP2$~�"ĕ���x5�^��yg ����dNڀ#�jUG��pcB����K`����6(!��C e��:�<n��\�6t�M��V:>��)���Y��k�榺;d
�~z��'-����;���Z��O��A��S�T�D�&��F�X�Ҳ���֧-��
���d�����**�|u/��o	����zT��7�RQ���j�ײz}�o�y�>Х�˶��� r�&!�ɬ]Y��	�6[w�� ��?iN��ڊ���z��ͺD�� ���#G}�͗�UG����y�[��E�y�/���sߪH����2��1�l���V���Ȟ?M�<��VhNC�̝1�;������PC�US%��S�i�j��w3����� ��( ���[��J\���OFO0�3��c���`��Y/�������AC��B����S0��]�(��7KNULڿ�>�U�l?-�{nZ�g%zv;XM�����]�����(����*���o�@ƀ����?��d9/��o]�~W��LEk]��(�%�Λj�'5ib�IiO����Pg�f�h˧ddY븝ˉ�i[�Q������q����G���Fz��16���߁��
�K��Ȯk�w�9U/~w@�XXJI�Oux8��g���� �eVg��4�$pvHA�?/�����i�����4���0W@���Zj{}Vj�V����sq������уW|)�`O �l�.to����dZ^�����[W�N�pe����?{R�n�>%N�$3"�J���Ҵ�)��c��A�#&%ZbjGU�H/k���U�x�Lg9L)=|��O�E(�i����V��t��%$oV&q���P���3�0��в�m��%bY�}e,8���.��S~.�%Y,T������Ao�K�&L�C�9L�ݣd���S�|TK�%�޸�9<���7M�8f�è4Ԁ�}�;���oyX���zCL �3�~�j�]#C�;Sm�H���:|DuCI@*�^�7�m78�m�����r.���+VH��� t��-�˦����>�,��gi����g��A	E}�qj���ҩpcl"�N#�Ks���s(0���P�dm��w3����f�`�t������/,5�f��o�2;��ʘ}��FI,�(oV�d$̈MeW�*�<C�Wˠ'%*P���_����u��Zb���g�
�L�t���?�P� ���WL����m���{c�]%��-n���5]�/�(nOѨf����d�oO�?#���,Ma�cque}E���a`��픣4W�ϲػ�C;y+�]z��<���z���94�p x�b �Mc9��~>uH�-D/����|hyv�l��f /� �5�^<Λّǿ�����F����x8�Z*|�E�!���"j2;���s����������~�ku������lHN.��0�{���4����)Y��C�!����9Ⱥ �`#t�/B�"��U3O,��]�ɰ�x!� vGkʕ���އ�שHǔo@Ke�ga���a'~*��Ě������7�#؇��'u/��W�:2�=������ă_<u(��c�>��'ypf�"$o������i���`!�_�{8ۚ�ԗ�v��dE�
�Y�@m+u�m����ͼi�����nm":d�Uz?s�e���Թt0�ҘD)�F�u3�#�4���[���\,�c�u�X�H��P*��`�����WƄ�w�6��n��,�7aY����tf�)}@xt���e
~_<�n�>u����{�~��BnyY=F[�f�[�=1OQёl49Qr�q����G�0J��Q�}�~z��`_{!/�ă*����47 u@�g��֠��؈�D�S��BcV���@W���剟 �}=��U�{�*�,A�V;�ց������+���O�]t�F�pFL�d:� �5uc w��&$�< ]Y/A�H@t�[
\}��B������h�~�=�1H=��Q/���V6���9�6Զ#�D5���z�ű�:VZw�R�Z������s1��.z"7UWa��F��)Cn���E���ϔ�Hp�j ���q:b���E~�?an��������8�LGB/M񧏺��ܦ��M�����ol�O.��cRR#����گ���)̤�,�tS1���W�u6��� ��]��&R�z���_�~�����)���)w�.����̴c�*j4V�g
�� �����f��Om�6g��E�,;�O�Z���� X��[^��7R���. �*�t_�c�#9Z���ԧ0p���+6���)��N�H�s ���c!A�O���~jM�BDά��r�	x���Qv�U�뭰�U���ڨ�A2�㫮lo�P�s7�g�Th����Xj|���Mh# -�"�?'��󍪾v�v�}k
~��~�懶�^F|���xYz2XC�!��o��u4�� ��o��u��u��|p���\�f���Z�~z|$����{�?�?p��"6k>X�����?>�ӺK���a����p?�~h�?\+>"�P�R�K�.U�y}���_����V�D����������,��h?J~E~(��s��շ��\+*��z��֏�$�L6>P1U�}��K}Z����w�
^�lJ_�����S�K2� ��e����Ty���|킩�L�9f��q�a�vi#z��*4�Q�����i���e���5��C?�-`�$��gL����A���w���q��p��Nl�P8#���;n����B	~wX�Pfm)�G<���6�Lx�E0���D�-��)��j�b/���UZY͞:/�������6^�XFCAz��&�Om��ε����D�aY�2����K΂�c^��=�I��{���K>�v��-.l\V@�bS��-��@���I���/m�?�.w
	 ��)�J�������$���8�/'�hsʪ���Vk�ƮCW]5��� ���ھx����X�-궉���}�K
�g�RSkܯ�M�$�5�r��Aa��1Z��/�
,�w� ���K��5�����_5�����9o&��LK=�g_�i��X�ᒶ��ӇQ�D�Mx��ޜ��-�^Ѯ�{�[��:�+c�U|�l�?]��?Up9Gm�����y�i�)�0N*���e6�cX�}G��7dF0�%�g-��ñ�vh	���>�\�׿������lv𻜖�!v~�*�S���\8$�T�0�����ս�Sm[E#sE:��N��&���u���m��{*I^o�ק��V�]|�tĞ�����5�7.�
��
DP�sG��R(&�<L�}p��&:�4���Dܮees��ݳ�"!���D�-������DR�{{��} �E'��R`�r^YT���V�l�Y`4�܅��a
?D�ȡ����l}O��)�����U�`�Mw����^_��B#l+4��u#Df�F����(��6�	v������\ԇ���p ����i�m7��sxXqʹ��{Dw����j�/�^�<L��j)e���Z��^i[�w ��uF����X��|��kZ>�.� ��i�Zx�߶A�} �� ��D���[I���xZ��u�V,V���@JI�^����=�y���O��� ;j�J��YS.:�->���@U,V�w���5g_C��Co��Q��4�װ��$߬Į�ٌ�G����b�،���6L7I;pD�Ξ�Se���/�z�`�l�l)�&қCmO2Ej ����l ���rњ����2߫q��/A��f�b�U^�a�>���|���z>�7�qr�TLm7�N]҄�@/�y�2\E?�'���I��v׷A+�$�M`�������*��]����@}l���/����l�j*��8N���b��^���0�p)k�sY
��ο�{����Y��zq���_�|q�h�Z��ϰ	}��l�?߳'��;��_�_�-�u�]ge�|����8[s�/� �3<b��s���PK   ��dX$7h�!  �!  /   images/c6364832-c854-438f-b38b-75bf2a0cd33f.png�!މPNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK   ��dX/yR�c  ^  /   images/d2af519c-c065-45b5-bffd-6bf239de2b90.png^��PNG

   IHDR   d   P   �	��   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��]	l��gw��c};��ΈU��ф#H�4�� �U�R����HU�V�z� �rD4��F��\���І�p8�Rb0�41���X������lf{vv����>�g��f�����������*�8ˏY&�d�xY���/�m\�BQ�6��#���a< )���������������~��f���rݟ���M�s���Ȳ���x= �IaB�� Zl�ۗ��������p�I���zV��ˊ������۷��v��/����,���$1�#L[ 	����t�ҥK���_����Y@NN�;wn�RRR�_s�â�Ͳ�e�[,>�7�AI�5DĐ�ˢ����I�&��2�M��	b���j����͇��cg��3,����r�x@c�0!W�\�[vG�p8���/���#�)��Qr��>��3L�9�e�OX6�FN�^(�1G����:joooHKK���"����.ܻ�e1�wYv��(�S/��t����P�������;D\I�Y��;,+YvRT���h�p�Ȼ�������Ғ3x�`b����M	��*�?�4�@�!�R�?x;��������/4A>��E�Yǲ�4W�{��(�ۉ	2n�8:~��~XŁ�Q��UWW�C��������Y^e��
&c�MFyy9�]��� e޼yqՏ�#)S��kg%���㏗s�=m���Ɋ+����
?o.?g3s��qLA��À�"V�k_�n]\�8�OI	���a��ڵk�9+2d9�N�&�|ʔ)t���)��@��<�zۇd)R�)���d�x���F�O��dgg��W2�T[[K���b�-�b�O�>B`�[�{������p�}RC&�6�gXo{�!��
b6o�L'N�S�N�p�]�}���Ni1w-�u ��ѣ�\�������h�ر4|�p��ʢ�S�Ү]���=�R��`8�)1���㡊�
�Ng�QSSC^�W([|���)4!H�"�T��u��bK�)wYY� %�� ���w������1		qdCo�B�p��R���L�'O�dXq;x�~��i6l�p�S���t����DEU#�)���y�2��SK��י �`\o���bU��1���@q� �Sc�����̌���A�Pt�K���7n�nJ�S ��Յb��[dS��o��f�q�V�Q��2(���]l}�4Q_?F�~l��=�������F���u8�)ܛ����R�2-�W�^d���is�uD�NXCC��5e6�u�LG+=9t�;؅����j������)/�y}����D�?蠃��G��M�L{��P�/�f�Iv[����-���p��N+�n A�&��y+')A�ج]J_�p�-�c\	N
̘1��/_N�������e��	VBA.�qd�̙��~I)h�v% [�Jo_�25ys�R���ug;=��h�����=[(1\���TO-���������tQ/+��2���Y�q,��!���l�U�������dy��V�WLt9����'��IA�0`�Ha�]�d	m߾�������`�cdn/��M�0!|��W�
f$�G�|���B�����a�r��.QN���E��S�e�l�t�(��9?�f�n$���,��4�jNO��"t$-�����A
Z<�pa�c�ܹsE9b\Z=������D2n��Ѱ���RЪ�����\A{/L�*�B߻<>l!�*զ)��qd�����.�a�7wO��n�f�=�<����nR'F���@�$��R��"�����/:yP<�-V�.�0ta �3���j-]����nѢ�lXHt�bq�C5����
�B�c�X݋Z|Y�V�T�����3�x� @]){��$�]`�� ��E"CF�v���`�޹�yp[pu�`�)�6�:�.�f����.�d@y(3[Ay�禋Q'��]U_	i�aAqA��ߣ�=�v~83"�{�V�,��1	]�p9P0������"�Bl!dVp] ���*�!��9���6_F�֔��Q�^�}(<�Z(�X'\n8}M��(
�Ҭ�4��2a!p;��mA�1z��gg �
��X#�fʰZ�Y�xϛ���1	ٸq#Z��髊1&��D�(n1&V�n��L�����Q���ƾUg�I��Ç�Q0��p�BJ��;!2�����X �C�Dn��ʕ+A�ZZZ�$J���28�T�y�f�}�>~ժUaRt%n0��TX�c<^!�,�IQ�u�����%�@�#�MT� ˈ�E'����6�=��z��B0�٤�H�L�w����!��	h����A���'�ǃ�	��SIH$�	뉢����!	��A�9�SS̰x�bw�@�u�������8����.��$���Y�9s����e˖)2�Jʃ>�zNN�M��֬"yܬHH�oD�F(�E�`�A[˒��e@�1;(1	n�[E�#�$����4���0xXPP�̟?_]�z���z%)2�?�p�\J�\��G��`���eI��X ����;��Z�;�x!ř� eŊ����ۡ[�СC�"p��c�xԨQʢE��M�6��d�HpV*^�q�UB?7�|������*���4�u$?PLՑ����<v��1hXb�q�̙1�����o�6��i)=�f�4к�:����yx?oڂ�0�����{����z<�=�-2#\�F�H�{���z	�~l����gY���O��h�uf0c�����>eVl}>�d��K�,ccU��P?z��k�Neǉ'�<�	E2vt����Ԏ��[�n5�V��$!�!:
����$B�/	I!��=ѧJY�"m9^,�!	Ijk{y��?��Kښa/��.*bJ�$$EX�tӫ���XxlK�dXb����t30��fڲs�ӣ�ZX�f	o�MZ/^ZH�C���늟���w�ÂD��&��$����38�MXXC��XK{5bU��O�諟It'0�T�vMu0Ȫ X����/�~¿"��t;LQ��'+}ݠ|>5�4��e?�v�߰%���?|饗���nX��,"-��;8��,{YvKBR��_+��wi.��1b�|IH
�ي��������_=�3�A��,��|��Q�\IH7C�)��+W�~��XO�e&��4ik�1�=����nF�UX�h�ol#�k��W�he�g����-$`��0���RFZF��F�e-���PW�`�ΨQ�^����>Â5��(�|6*<,	I�m�ǌ�>��e�|������,��V����ǉ�H�B���z�����_��V�B�0�.�|�4��$|��9IH
�q!n|���k�}bj�UB���9�X��]g�0�����V	��=�Y��D"��Κ�7�,dYb�|����$)�d@wm�����0)O��)B��fA���u�u��l��"��`���N���x�]?�~���&�e�_w:�x�$$�|��#G�|�ԩSq������A8c    IEND�B`�PK   ��dX�'k�  �  /   images/e8452abc-1b33-4025-a556-b46ce3c60df1.png��PNG

   IHDR   d   &   2r>3   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��[	�U��j{���zI��t0i�D���H$��3g<zt	G��AFe���(*3"�":.�
!,*[�$d![�ٺ�I��o����ߪ��@:�%��Mn���������zo��{r:�P$�����Jv�W��!�6Uuį��뚃�I�Op~�/���$�v�a�Pw��6�>j/��n���G�6�Tt��}l�St��~�S�J8���'����ċcÊ��h:��<���c�$�	�4@��}WM-M;0��Ј(��n�D�:��朵$��x���D����!G��t?���k�~�����]r��4�4��5��&E�NxO��i��}��\<�a&�9B�o�؈Ӹ�>�3+��ry�]T���C�ُ�ˏ@J�ìkA�e��(�϶��Έhϵ��3!��ܹ�!U�Ba�]�p!M�͜�'�Po!�8�I��sm���}瘊K��de��`?Sk�����^����i��P�"���b���LD�	��0/��ٔ��LB��:~b��*4��t����9�ae��"�K)Lȸ��t�y�GE[�e�I�Nc�W~d�⿎L}�B䉯���\a�d��V���5lL��1P]8
&]h$~�]�,��D���Wqd���t�p����1��jS�_[!b�tϣ X��B���cR�Z`�<X����2Ix��<ԧ,B�$1g�x��qV�.^��H������'N��B>�X�Dm}Y�ܰ�w�G�'f�y��h�2�r9H�	��gM��[�K_�aȧ��R�	է�fT(H��4 �^�&��P�j(Z
REx6TG�9LL1�z�RqZz4��A��"���jנ�	�W��U.P��m�ϩ��% W���ʑC�,&�� ��n#�D�j�Y��r�n����{�}�,`�@�f��I�|#̴i-T3n\>��щ�΀E�i�w$��� fϞ�k�����'.f���2A��A���~F0�'oCJ���(�Ť����j�Ѯ���h�v2�A�tt7��ۢ5I�+��>���� l^�;mC���v
%Ocڇ�N�!=z%�1���DL�����S�v���(�l�EA*�&��{;��ͨ8�MN:1t��P
�;��D� �?C�Waeft�Ǖ4�E��cČx@#f88�ȣ�&���iHU�h?�O?�$�.\H�I��4�2\��p` �H9�~�s;��/����a����0SK�*�a}V�g�F��b����&b�Al���j���A���o���	�]���VPtG�_~Ӆ�k�m���Q��`�ԃ�R��k����ކl�h���|F�5�����=�8O7����G�M����.�@�������G��Ryt&Iw؄h$	��":�%�>�Ïko��h�Q�1��H]y;ꪪn���K�޽�q0��Uo�`�RF����V�H�J�O�IT���Q�OP���$��"�
�L�k)/۵�8��6�I`ŭ�G����q8w��;y�y�������0=��D^��C��/K.,��E���4�T	�����]�<u�.���!��XJ��������7L̲ϙ�2����/���3���Y���1�"�L���%?_؞S&`�'��z�ʛl����9q,�"�d|�T	ӟ��4>��@���z�ۻ�%��!�m�w�Hr��A���+��@:�����A|���&�g����_��IÞ���u�1�y]���e�#PN"!�Q=�?��*b��;���j��i��Sf�R���F���,�aS0l��q��ڎ")(ɒ).��֧���p�Dmď�����t�CUdl>�Ep����i��5k��U��/�sd0��cv}�����m��xlk~E�wT��!̌A;�����R�o�pѠ�|-�WJ�xӨƄ�$:���H��X ym�E�R@��"����k$�:s y����1��fƺ]�8�>&^k�ϒ�G�X+�j���}�\��1�9g�^�eTo�z�`��}fnH������[qo�u���7&p��,_�4!E!�@���-˂��0MS<�w��4���4#&�>g�ْL1��]d35W"G��5̫���v�k*���֭_�K�/G�$���(b�`��T^����ά��C�;C�R�׆��Л"�9�Ag&���B��d�������4MS!Z]�444�
݋��ATWWc�̙hmmEKK��$:::��da|r��Wa�Q(`�h��Z��[�$DolCb������"�Yd�.��PY7�v*++a��0�����Khj�~�k�-|{;��e1C2��!L�

�V�x�Ј#VD0��e�SIn���V���)��kjj�`��Fz��؈T*�={���`�����*��ӧOǆ#q����c�k����y�SEL�H]&�%�m�=C͋������'��ޡ!��ރ��[a�*q�3����%��U����i��r</���l�\�.�ڱ
�)*&�E�ߧɱ:b5��:�Ţ`��g���+W
	:t������/b���طo���3Y\gFB-Y��&���M�@��*�dڞ>pS8�HӸ��B���a�����+?F�#�@	�g��N? 
&���h�˒</�k�M�;�I�ò��Ff!6Oɴ�
�^�7n��ȑ#BE]v�eصkv�܉ٳgU�u�Vq��ö�L[&~%<�� �-%�7�I"��Y��
I��
RY��W![�`���~�0�n���/aْ%�����˪��W���"����'�"�����F����Q�|j���N��Z�C���ǠdNڊ0CX-����Lٿ��f�Ē��mmm�%����=y�5Va����TY *Ո�
�j?yTgTI9�.�>2��:��[!�Ůh9��9�%��S�e-�z3�;<�� ���ݨ�6�*�Y �J���͛�x<���.tww�w�Vx��ѯ������8�3|4�O`*���0� �xW'�ɡfV�D�qp ���]��KR���6m:ló��a��������J�A��]/���"�ߎm c6��1���3��[UU%ο��jkk�!����bH$B���L{Y\�Btb�b�؅̈����	l��p2��$��E��� ��]���[��d%2��E���Q[Uq�/�o.�UV��@-_0����w�<<Sh&�0���l?]ac�c�aJd�ذ�
c;�##W�=X���0q�3���H�H*~��p�]����ds"�ۆV��ae�b [Q:k!�W}�?܃�tF��H_rl9���L���{�xte݄w�F�xU'��J�H�H8n�$�P��]��e�a/�$�y��R�2
KP]��Ϲ��zT$��y����Z�.���B!�-"g��/=$vk������G���éK9!�(/�=OpM�-��:VaO���,I�>	/�\Ċ��w�Q�Q��R��Ҕt���έ�A.o_�("���_{����}��f�~UxY%o?Čס>�?�{�~Z/���q��[��!��ea�Y�k��7L�QJd[.ֻpsh7μy����E��f(}�1¦,$r%�0�"�sk�¸�����J�w���.���_}��H]/k��4��T׌�6��؏.+�K��g����'��#��c���y�`{ ?�R�_T��X$5ў�(�.��l�Ķ�j�^�C[_��T=�����5/\��������tF}Rz��^� ������G���<E���L6V�L�퓧������;}-^'f�j�Ϛ �����EBIlPu�d�He�����8�)�𲊤�T�!�����?q�w ���#b�4�}b?$������p�|Z�P����8ht������K�N�ca���$�r�֏���<�t��,bjysJ<#��k8r�LT�,�h���y�}���Q,oCJ�_>4a{G�n [Qj�;�V�A�{�&�
U#���Zɡ\�����ק�e��gޫ�]C#�a�E���ӝi䟸��xj��` U<=b�;��7��[����f��:-���D�������8���i�i������.���7�v�rkx'��y�	xp�e=7	/��H}��I�v#u���҈؆��_T�lV�8���b/�S��i�dJ�ѕB`�;E|���t�b�e�q|Au�b�w0��f�3T��e$��׬���c΋#�s�nO������%�І^����\�d{!��Mqa�_h��u����"�4U�9�B)ً��F\r�%�'��
��kXa�&0�OQ]Hu�H.�=�c�əʹ�*���O���"����u����1(�%�"ͺ�3!�&�� ��V�~�Ex]i[��i.�[_���ދ�+V`��,�C��s0w��7�r�8O.2QC�	��/k��/�,sl���-�.X��Mq3�
�K�HNID�?�^>8(��_U����3�\9H�D��k��{�݇������-!�`(�_�����.��D�����J*k�)TV�038U���������,�����Nz۽�%�G���f�7�D��؉eq"��� ��N�6g{�,�Y#�!�Oo�}�ń�Kj��a��hy��]E#��}�uw�c�j[���_ �ę�4T�\�=uB�M8>l(5��%�&v�!�:�?�;�fy[Z�3�%�ENw�?�ݬ.80s�|���{~/G�!�a�����
Q��;q����#��A2�<�1Ln��a����,�8�p�p`J&���?��B�``�t]߲C'��v�Z�>D����ؒv�~X/ݏ�?܁���U������xO.�b��)J5ᛄ�§6>(����	o�q|�y�J��~��(8VKK���و�l,F3��S���.��	}��, ,i|�y��y��!�N�sv�z�"�N��&��k���l���a���z��#gaQ�ii� ���K�����6ࠀ�IZ!�#�l?����1��L�$�RQ��qR>>�ʛ#g�X���:1�[��&>�j��Hö�h~
2�e%&�e����P)��u�Øla���1#*�8gh&��
�wh}�P$Q��SDJݫ��d�"$	�f�CM�6(���K(�"�22�
��W@%��I�p#��C��E���-�?(#�Ȟ'ٌ����.t����)��B&<Z��:�'=~��Y��.�U�3�����!�P��yc�/�o/�]�����������I�nTV�q�G>5{�������pw׎HȤ�����>gP.V@|` ��r�	�L�0����2��~K�+R��"hOj5�U<X��dZ��O�L���:n�Bm��d�'��T�{��M铿I1�6[��`sp� f�DB�%��/#N�����a!1n!E��`��ջc=�q�}�����d��\���yMu�&�eq>kX-w2��b̟��HB�I����f��ؓ�ėV�G8R��FVF{�5�{r2"�#v�
�9��mT�H
�̔B��}ҲX�C��I�o��ICn�N8�.#k��;�2>�����6��Ǳ�`�!i˅� �]��f��q�](o��G����9�e��:Ё�S��*��b�|d��E���םX������)�؋)YT.<�<Mܻ�۽�M�W	�I�h�{�X�3��wƻ9#cS�]F|��w*�������������G������ß��go=<��c���79Gu�T�iT?�';T��G���Cf/�jJ�A&�	X������KD��'�o�
2�Iˆ��    IEND�B`�PK   ��dX�+�s;  z;  /   images/f3037bb0-f56a-43e4-a2ff-17056f7c669b.pngz;�ĉPNG

   IHDR   d   d   p�T   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  ;IDATx��}�dU����z�B��=��ff��a� E��~���bXu]W�[]W�.:,b �H�!ϐ����=�=�su����ι�UuU�V�ou�Ztͭ���{���p�S^i���6���-��d~���q����n�%�c)E�Q��m2i�΅��Xi2S,��'m��.�FQ���-���Tm�����b0s�;B�~����e�>'Ax���;hW��������߾Om�P�-����sC�z�C�"�"�ZȐ4]PR
��m����5�������(|��D�>u�
e�ڶi2O]�m��$��0���9@m�������+��XҰд�OP�1,�|��� ��r�:�P�����:駙9E�)�3��5Pn�H��~{����mַ_��|���O[�)�٩����~qme����
`q���eIm�ō��!-o��/@Zє��7�dڶ}�|���m�
��-��!��he��x��u��6�o��~������_�$�.Z|��/LW����yf�!������o���h}/�|s�o5$��`qQ�)^�Z�,�̲��n�V4��8Ǧ=�`���e��J4#f4���`ZNѵ�iM4�h�Ry@��Y��3XL��Ч-F�����k6���,��LW���a:U��!�����
�<�.�0�x��N詔<�Q.�f�dw@���H�t5�C?z�v�f�ॕ�g(x����sYRa��]�^��Π�)�Ѡ�fF�Y�o0��C0��+p!�h�Iv;�H�8]���՗
 ڟ��h�4#��H���A<v����A2ɫe�{��caV(�(�Qiy����X����3�W3��@X��?�EI4c��j!]�"�� ,d}�D׮[涯�xSԥ
�3�2�b.CZrbe,�2i#;}Ƞ6�d5k��x�X�F�`��h�o\i:㼹�o�K/<��4�Mc6�*�Y1�g�b�)�L��E��>y�يܺ�652�=/�P�mWHa���H� M��Z
3�3B�����h'K*Mk1\��cC(?z of���.j�X�d�X/�Y�Ҽ���n��iE���1kD�͊��u'�_Q���n8��c�n0e��ym�à]2��ߊ�T�u��=��,�~O;�;=�K�n�"V�G�VB�zR��GV��D�q�[�Y��[.-n���Y� M���1�%B��Y�R3���������Ĳ&X)��X�X)\N���8��������{~���*��X��4#��j藃B�dY֓�P�6�t�H�����f�̥��>�Į�M<�U?!���|�}˜϶ؙ��<�����6��p҂���nz(CT��>���]���߲����[�D�چD".�a�.�߇v3"�8!iU��[ݼ��4j�9����#�x귏����c�觕o,}~�1��WRʂ܈�4�m���$/Ȑ1�6�������ӏ?��J1ޱ��,�u"1":���L��qO�Ik�Ѯ�!:�PuY1��+#1T66b� �x��)�E�z��P���ebJ�p!�BMQY5�=�@_��y����s1��҃ŭ��՚-�]��}��`�Lc�4�E1�8�hV҇6{F�+aAMezN��J�Lo�$�]]���u%P3,�)�c�D&����&�������D��ٝV�J���54���[`�B��2f�V;m-k5�uz0�?.�d��8M3ᯮ��ӅvR��OΨ�l^����C�3���'�(�Hf��,�o�&�^�n�^y�;_�n5m��F<���*�d�[�8��z`��J�`_��D��;��!��VRן,s���@g��p8PQQ!��O��eg�����)Y(��;��o�.X����ΚfX��0x	����k]#�k!;w#�3�:넥PK�C�`���:�E���=S\\�?���H*�Z���Ls�K&��H�h%h]ؾ�!<���(00�L*-�|1q50	}�82� ���X�N����o~�
�;C��W��";f�A�Ě�O���P�a�>2u�R*QP�c+t{0��|r(�F����f�ʈ�g6�^3܇�ۿV[�\d)n���e������Շ�o�C~4�r��U$���i�%I�T���좉�!��:aŮ#�#��Q�%e�����E���}Q�����<�h����4GؿEE"qv�ˎ3��B �%s�%�/- �3s��lᕖ`+�f=+��i�\f����P�I�ξ6}��-v~:����-�CH�&�|���{&Q�b%�z{�EgY�:����:������m�ɫ:��x�x�w�'���]�ǡ�*�t|�܍k�����F�UR`��K<��[0����o��zW�>QgGR�����'ahC�=�ъZ����Qd"���z��ƞy	�?7	�Q2��C&6������ߠ��sz�p����.���HX�2q~>����Iv�2ы�Ƣ/�'��g��iH�;}U�V�
��t�H��)�����0r3C�0������$��̶<p)�m�o�9hi�HN0>{Y�����E��CB�i|��jH6R}'�����4A�kj�*L���V^)�(��a���O��@�k٢�$��5@'"9������D°R{=Grt �8�d��Zh�{��TYEmbЏ����*�4�3�K�ӥzV�Ok_h�� �B�A�C�n��g�gƆ�coB��Y�����j�7�L�����	�W�L�c�]O���m�.[����u��P򳏣���a)��؝�G���!����|U�y��ct��H�1$b���gP���g2��?���J�$������-����v���'�p=���^��@/��%p�{���;܏�+އT�a��䋯��Ӆ���,�u�QMe]���G����:
^�!=Ǡ���#���,�C�����X�H�UP�e�p����lM`5w�.\.�f
7N:;(�*e�I��I#�JqzR�}�t��S��B�ij�V�DM�O�����]�@�O�~S�Q�-�
_K�*�O��Y/�Eu�?�pԏ�6�c1�%��t�sa<�l)�bvH�woC�?��.+��4�.�i�ҎE�J�5��@Z���"�=��Ϡ�̷kl4�IHU.���v��t�LP^�R� �i�T����5H�hB�:!���	!XH�����-��ό�BO&��0��#6��C���T����a�R����Ӣ��	Ȓ�>Mb��!{�P��nc�)�,>3$2��i�fxኘ�0(Ғ:Ns;q��C!��yU���S�c�7����k"@3 ��4�ii3S�y�Nz�J�X��e	v�"`�;���:�B��
A0-A��;��7"��FJ��H�B%]1y�� ��Ĩ(\OO�c�G���DL��J�[�x&�M0I�F�X�'��oC���n�`�D��L���H��hZ��	�}$@D�т�1��y����|4J$#~��I%��f�"ZS��� >�>��UM����f����v�_Nm��5<��`�D�'�UX���H��~*�#�l��*����C�o<uJ!fRC��0�K�����Y���ob�F����cV��?�=�x��&��e�~��%=
3#��U^�:���ue�8�)"��9�"��b\�~9��������i����7�?D�_nw��M�L/��M��s���s��9;d�P�=�O8V-2Z�du/FN ��_/�ȱ!�0՞v��}���%Bm��ϬϨ�0�zF�N��GF7��r�i[8](�X��uE�������$�����O~�n9c7]������Ӷ#��au�浈%�L�o�Z�E�$&�7�N�Y][��HN[��� 95�W_��	��c,>�N��w�����n�yYhln�燈����k���Mm��a�/&�Y�q=�B�lFt��z�G���0�g��9�^���f��� �iaC����!۬8���9h��=p8��$@�
��h��K������o����VU��uo�R��[i)DШ��d"���
�k4{�f����@����Ց4	�z��ڲ�O�'�E@����MŨM�\�v���k�ꢬ��xt0���T�(!�p�ظ}��CH�;�g�����,����K���Yh���!�ӱ��t� �L"M%�CX�*o>�?��C�y�dt6�����ק����g����eE�>-���/������x�p$f�8����ԑ� ���Ț�!�+��	��ʜv�=Dv����N�|�KA���7�B�1)�ljNQ}�=��;d�!�H���3��=���@s$�K�feD�f�C$FL/ll��;����V�<��7#�XN2�˕v2jB�˝�@�����D��k:��߷dt=Nl�p��\�5&�tQ%{|S��3C�sP� Ms�Éd<1�������d,mY��7�wS�_�wi�w�4��~�~0������Oi�Y4L���%�00HD�&R�F;�s�"����*��;�}���e����v���'F����f�&�_}��}�:�Ēp��������n�IcwN���:�r2����l=��X�픭��２�����׊>؅�������쇢1d����1r�LzA#���(�"�P�u�[�!,���сa������rܰe�	?��r�B;�Ey��a9�t�cU�;ػހ�؎��!A#�$��meY��s�5@����2$�	bH�]2�t�1c����\=�	v�����;��=32$�}n��a��ײ��}q�"��8��
�{��@������1V��@�4'8Dk���o���",;��-ȹz�����:�A~��ާ龳�!|����v�a�/ːI٭�myF�$��bV����b��w����A1CF3Sǿ����
s�'��?%|O�Oe*?v��fq��e3����-4���F{���>���^�f�_�������2�nN&S��=��b�,1�E�����F�B��b��n�Ӥ/��a���r�v�z&^Vp2\�2�'Ơ%�0Ek���ԊL$�����Y��U�����@g�^���#�u��{��뀕���2�#ƭ,J�}Ub�����R�B�׳�a��HRȯ��"���J���$�����
C_�sti��2-9$�)��UX��k��D��vH�D�}��C�"r
e�\���F�H�����.F���_q5��
��m@��qq��K�@���&�x2g��E��h�_��I�\04W)�Vݢ��(�{(�� �~qY��y�~�5(�{ 0=��`��P���pd4��ë��ِrb�x�LJ��W�vHn��gZ���Đ�e5,En��ȁ��\�$¿���h�I�7�#nm?�e�����]t����!�~z?�'3��hVL��(+�'�'�![&�Q�����PgL�f��~��AKP�@.f�Ёي6[��\�~Y��� ��K��ٞ"�'q�z����Bv:Qt�F���?���W��l%2�\3�r*��������)l�횋��&
�b�|6��٢������I�e2��8�W�2)5�XA.dk�������0���,>�\�[�b�W�@:�l�Ӫ�8�!C�.��]P|%P#!�D0�³(�~�����
{0�QKƌQҴI_�@xYhN4�0��� �(%�BɆ�z��"Y��j\ͫ���#��+p4��:�t��u#?���V��?�A��v��(m���b���#(��5��p��'VW��?$¶��8����Dp��g!�櫰U׊	ȓ�VY%Dw��A�ܙ0� ����m�VQE�"7��ar��L�@WS�@FB�Zb$$Y�s��1A�Ǎ�l�8w޿�E37N�1	 �z�D���C��XfxXYXD�XQ��fأ��Ӌ������G&M���`	b�ٽ��	�[��i'��:Խ�dB�GM��ޤ6g	z�{�i��썶��iO�<t@(��Ѐ�<�N#������V�
���;���$���[X:�z�ɈP��(�w͜La1�Ngo#�#@���pVz�a�Y��ٵ���2�cN�هk7��F��wb����U����H��B+�1�� �1%�oG���D�o�V��.�/��s�a�0_�
�e���3�Z����d��ayE3"yi�y�V��AݎǬn4�^��[����E�"�cq?~/��2:;;c�_V���w�Ia��~<m��Q|݇�#�X>�vZ��|�k_�/cC��=�1�G�B7�T,��A��r(ⓗ�gl�ǯ�n�:&,Di#��L�W�G�n���?�{�)���"Z �a�i��amA����Ah4I���'�4��p䅃�R�(�P,L�J�*�|�g�A<V�̄��-�i),�憢-`e��f������^�+.�^"\6��g������><�������L�1�q��V=����i��W�{��N�����&Y]L���$2v��D�B����C��'�Z�] ��
;Rezv�W��-H?|nR��6!nu�%{�T8��=�뗠{Z!�H@=F��ƿ��+�<�V5��	�3*I�S<�[u��ۧ݊+;����DҒ�2�� �ǘ�@~G1�~��P�?���9Kt8S1�w���x�[��~��⋌|�drF[�ۍ�r����b�)fw	�X�f�Kb,��C���aܶE��c/l�r��c>�b����!��C�¦�{�|��HZ�yb��V��p�57N#}L+��9,��}R'��>$��ܷ�����k�M������ʍh��M��'0�ė���-���3O}�8�u�pa8�"1�����%m�`.�p=3���'oڄ"~�9h�h�ӆ�n���>M�L�q�	����$��_R!]��5lw([�>4��<#'�K���6v�JvY�hʆ��
��꩘^6��>J����U��'�)�$%Oޓ"�y�Wx`�bC�V��eZ9�2��-�W^u��\�(Y@��сM��b�E��х�9�f��!M�C����ڇ����a�V�qZ���c�A8�[HIy��@�	B�_�S^J�,C3K�Y�E+��bS eǓm/f�*$�����6��d;_l�r] y!��?!�0����g�M��9�4pk;w ��DG�+~���tE#}�o��+j��	�� �(p�%^C�=.�Sߘ<�@�Y7Ŕߡh�W�ؐ���%
B_��͹�"[�Ղ��}E4�{C|���p�Q�dВ1X\ޜ��=�(j�:�&�XYY)`��~���	/��"�2CfIr���`E� ���F��w���;9����p(�7P7N��,%���ɺ��pVT�}�K-�U�\�>��Ŝ���0;6	�{��%dx}��_b�m/�ɑc�����,8�>I�e���R#1����*w�\(++CMu�	j��̙���ƻW�p�d�$�h�����'�R(�x�ڍ� a�A�rF����ņ���`�ß�{��<�JL�~�= _x"0�
N"�ԣ�#_DQ8���/��D�\9�+#!�]�E�2��.��d���
��p8��H���c�/ Or�I[,EQ���x�C�#�#�%��=�Xk��bt�0c������5t�n�v䈱`��K0U��g&̸'��tc�3��D��|����(��:Ay$�e��хzlJ+�EO���a�H�����pCQ,S[60�i@D�0Y�G��!f��8󯺺5U����#����h����Ç�q��֬�v1��*2��xb���21&���o3�~�, ���֞��}�8�2+�زb/J<L�4<<Hv��N��*n�?X��"�,p��!UUU���LQ$=I�B]�BkɴL�k�	��-R'(��D"�λ�����+�PRչ���l�%.�,���B3���hoG�"C�|[+�o-��V�sX���&e0���{:�%��԰̜?3z�V�ɑQ\�e+"�Q2��ˮ�h_m�ˠ0[U#G��{��̲"]ŵ��7^Ƿ�������[��pS�EL���FaUk�1����ۈ��|I@� [�Ծ��ń�M���[n)@YYg�0������,1��Ċ�8ғC`��۲
�S����E:�B�Dn'��GM3�FY4.�ˍ�d���Uը��Ĭ8���	�&�U���f��b�J7?���d�󷏡`7\֮]+c�I����}xf�s(&��,�l��l�㍞�4�5��e���@g�S"��}Y�#X��0���(��*����`���;	�T��d.I��4��@� ��P��]������8����F�57>�������>E�8�����Lx���!�Z�
M�a=�H�����µRc�#u�PS4�Uh�i-z������/��T���F��~�`��b�ϋ4d`` c��|�=Z׬1|\s0�Y�q�Dx�wX-� A���7�N�I���	T�!�h&O�m��+�*��[s)uj;��Иe�p�Y%%�������8�����~�H@�0S��q>��=�^{F��`k��\B bU�z�n����@U]����
l�Q�����"�W*.���D�*u����&h��D�z���3W��4F:�	x�⢘|ԟe�n����*�X%iى�{�xz8G�*HӺ��j�n���2�/L�"�Yb���8�&�M/̈��^�S�I[�I���ҁ�"SXI��e�S3F:�}�#���	|M9M�O{��]��4S�؞K�еե��|~���9��4�	�zpa�	����:��'�Q�NzM���l������.f�[IR�$�.�����!�zc^��Z�
Ȭ��ŃH��%f�[Ҁ6��Z"^��Ļ�}�S�np�EƲL7��PL6�H&�Ԝn�̭��s��%9����"�W"�����>�n�B�m�&l�&��<Y%�c��/��ƅ$}�<76���ǡ�3��7�� �Ua�I�����~�N6��[�R��a�<�^	��):�O��}8j+B�KAM���(F�:�*m9^�n'n�����p�ھ����Ӄ&E���2�W#zp�'���ߋ��h��ۍ`�	|��# ?��ag�x��Fr'!\'G�n>�p�x��L�-
��FFFP�~-���j�oWz!�IhW0~��aTUV���6��MU��?���M�Aó����7X�В��t�3���>�I��`�-��a��j���c�h.;����a�:Y��e�Wxx?�������=d�0�a8���|�)A�އ{t'A͙��YtG��Q�i"
;;N��|@A�P&��:E�IG�<St�2��|4>��b:A�k@(�0��DC��**��r/!}�z��ć�,Q����O�O���&K}�=��1?�)��p�s������y�#�8A+㹗;e�w;Ĕ���G04�4 Y͹]�*xq��Z��>.ғ\�Z=|P�K�rx9��l�_ºj%��<���ݹ�!|E�D���"��Jp�����&{g��{��9��� w[{��}��dk:�O�'��
�A���A�P19�uB��đ+pP��JJJP[[+���ȉ�jG�E6�<��|���R���&�1*�d����OJ�.H�z�
]$�͟��̨&��!�:Ja8hL~�����;}�L~?�L��3�!��8qa�'w�Y6��#�����_Ax�F��4�������L4�e�턪&V��k��N����Alڸ�_v�ܱ�>�(���66`���@��.�9b�X}%�^?��W�QRQm�(
�$<�.!㩟�ub�h*���j�e���+���#�����\e�����E"�|�>LsJ�M�c/��.,��`I���C�xP�_�au"�X<dHB3�Kl#�"�;���՝��34�Pz9M�Ёɭ�D��Kn�-[�o����.l�$�b����[�ك�^Z���G��P�����=�z��`��M��T�JZ����N$o5:6�[O���}b_���+Ѵ��h�x�U�2����=e;��,�d�`Ög���[C��~�$I݆h �FZ�	}3y�\YfH�~��L��$N�<�#�w=�����Σ����w�p�͂<�椩�oooǦ�N��%�}��b�5]�ޯ�iSv�p=�ů�g�^{�G��}�qU�r,�4�e�d6C��T��6�uB������'D���&�E6���14�M�P�#�1��*���g����fiqĐ�-�səL�����	#���iF�S6�['tF2�p9{���c�Qݼr�V���C���x&����g�_��ݮ���\�"T3��=b�o�8˫q4���چP,�DA�a�l4�W+	\alR��#d9��������:>t@���"�Y٧zc7���jY���Qw�����8����w
Ĕ�;Q���Rz�%����V��N�(Ny��{�J�uv��!v�gl�"�w2��+?���"�/kF�nZF��>�Bg��\�ؽ�m'��ϻ�x�`�F����� j�����
�9=ة{jjs��J7-�GFe@1^8A-i�1x_��&�1-��3�5�l=KlSQL>�4<��F�����M$F,(jY�T_����G2)n�8�H��@O���#�ۀ�@|g���+ϋ�
����!nK�Y&E޸|�����>�gt����Ҟ�獻�%��J��)���g���:Z��Hϓ�i#��X��o�.i�Wu<��,������蓄�톯_2��L���[$sv�M:jz*0�\�;׵""�<>��\,E�[o�,� C=��C����aD��`�!��@"��BǏ�H�y"P7���u?�G��pM ��S�˼�e���Fq�v.Ab�cɮ.���n#��!+���6\�!�^���$&�T1ƤQ�;t�C��=C4=��+���QxRQaq�R�s���=�:'iZ���[�l�d섽�A������u(�����dMK��J2�q�1b^�9����Ȟ�#�W����Қ�:q�
�q��%��O$MM�ά��i���x� ���	z�]n��WP�U���v$����b��P �w���%w<�˗§�IZ(�+T.ݶ��v}��O��b��^MR"J�]�+क�	؊��4{ݰON�E2:v�؎�&��(�B�f�N�׹�T�[OB���H���-kB�d��\�lTo1ĥ��2MԨ��1�Mے͓���0c�o~9p� .��,�P�n$��;O822��=>�.���J�:W�3!r`/�$�#���ZS�T$*�a:[�����!��4�Oı1��/�U�\���~��.x��Ι����v�vثV������?*�Qݼ =|5�����q�kP^���ŞF5F�՗s�#���{ϫ�QG��b�J�J��-^�3���J������*D{���E��R\����)	fV<����N������b�����"$߽[����w�}~�[σ�3���?������>�?R҄�n����)���	f����[�
S,���'1�%��r��r��mr�K<��r�6�S�y���c� 4;$�8X�<��� 0&i���?Ɨ��c��|���ouu��F�ܫp��X�Q���h"�,��+���z߻Cl�)�~´J�6��!!N����9
�(Ь����8c����/�燂�V��Õ��V�E�
����bqó�\A\�j���&�����w�,2��kk���l����ϣ%�%`�d��0�����!>�����y��D'�����w���s��>���p:��M����[��Zojj��3�YGɱ�����[k)�+�ov����Q>6������4����غ��<��X���-JHS'�H����Ŝ5<uޡ.�ϲ`�D;���`ǵ�@��Ni������POn�c~"C�H�ߣ-�{xX�>��?���ċ�}%#����
��8V�g�Y��8�ÿƱ�n|���ओNY�<Ax�d0�ǟ~/��Cv�W�ܣ͒�Ęs��/}5�ӳ;�����5��[��}��nNv��F'o��ྀ̽s�y���H�Q�;=����[}����H)(���o5�!��J��H�1�ɨ�Bh���0"�Bm_%��co�����W�2
�3�g����뱬��'wubt2A"vj�q���"S�"�p������GCC�4�]�������H�h�T%��&5Ǵ�[�DL�N�\V��V��kO�ˌC�/��T��N�J.��.��|1���nCI篰�p�8�)CW���KkE�n!���`�-��Ѩ084�~���wC�"]B�L���g�j��z�2�#�ܗ)ű�w@"�u*�0���7� ����2�f��ĔS��X�j� ��{L��s-湓�D4��]9�jxz�{F0H�т$=��컛&�
p{��Đ�׈�-�rbf�<x�o�ג�'S�֪
�%xxx�ؕ~୅�>H@`�.>���"�S���Hv���a��˅b�/3؉u��u�p�}⁹�����ԥ��V��Hb�}�rk������$#AB���1O5�����n!)Kbq��xN^�Yc0_�����Z*�X���l�t��!��.���^ ����rb�˛��ݐV4s���,^���&^��o=.H�{HR�y�Z��� ���9�u�J7�у��Z�hʐ��م�"ZeV���4�d`n�Ԍ5��3b�F��S��S�� ��E*?G���P������˦��=4�Q�ԧ�:D�w������01/.[�=0:�	������II�e����i!>�ה���5��$�1E3�2��դ�V\',vf}=��+�C]���!5��!J��o����^%^��o�.|}7�)%�'�@�h:�}�=��P�~9;��_A��ԋ[x�X"�X�J�����I!9����O[����@H��,����Ѹ�L$11a����,����pd҄G��IBN���"@F*G�,�XWg�{(,��܌6�y�t���Z-	�$�+��_�u]����Q��J�af�n�b�rb����Kj���̯�f��9V�"� ����@?�À֚��Nf$�)��03Z�u���{8���&ie�=D��_��H�S��Ey�6fF���A��/6�#qw�/g������z���p�l�ĺ�:���rPkYC�@asÝ�Ƥd�hξ`�7CK���O����<j�A2��Vd72�x�&o���k˪�%h�U�S���4.�[`#��&�z��T���*¦�H�z��[@c�j<.�pXr�}�b,	��������mB)zV��.�D��{Ǆ(.�C%=8��Wn9y-�����`Z�����eZ���gosh��R�MZ��!ۀ7�Z��;�$⪞J䗳kO�f����]QPJ��C𰴴T���WI��'�$���Cq+�	11øp�>��9�<���J�-ƓP]�VA�ׂ��W�U�}N�Q'�l�h�NXeS.��"��yC�@Y�?ہq\��f?�z������ET1�.o;k1Ђ�>CY5Ը�W�;V�-�O�<F�W�31�ҿh�2����}�����w��V��Ob��^�$��I7�����Dk��ܲn��د�DVn��n���K8W�&���w�Wހ�<⽯55�Ѽn\�R�߭��O+���B(k��k���r�D�-����)B5Y���G�[i���z�O߄3�p1ڡ����E�YMm%�VTQ8b����X�B*�� ;����I����,�Be^�'z�i����l����al�#��<�.흃�b����q����
�r(�t2t�3���Ca%[G�ض}ݍ��
.!yG�u=#�]����~X)��l��.o�U׊�B�3��S�.e�H�Npr��A��$�O�/Oo�K���P���	G���=�����xd2��[��U)A����C�2��e\���À3������$z��X�:q��d�P^b��t� ��G�f���V"�d��#�ә�+ԔP�)o����K���7�k�"�A��~�zACS���$ho�3�q���.~��KjX~/M��km�E�pޣwuؤ��c�W�V\0u��� ��IؿV>��V��SCp�+��2ـ�᰺G���BmGt�V���ŧ�,��&nk/rQۍh?8�J��S8�����ʋ�9m�� ���D�~"�l��E�E,�~R�c�e�H�ץ�Շ,�ʺ<4B�.#��M��&ɻI�3����Z���v�b�b�c$	4e�eR���5��}�m���~6Ĕ���^�i_���O��Ж��fb�&7y����c�g��$z�Ľ�ޏz��`����#�ȐcCLl�5N���ࣻ����bbV1��Lz��ڲ@R��3�1s[��m9�C�k+e?Sǜۈp�OL"�A"vS��2u�ܘ�D:� ���|.$��䤱?�&�B�L��mMNX/6��2F��ߊ����@5ι/���Ǡ�qz�S`9S�C D;FS���z��&fӜi?��|�-��?�
��m.BUg�h��AB�˃=�q�]x�tG��T�����q�\�I���e��c�i�xz�lgP��|���ݫ������� ��D��s�F��>z�7��Czl����`�&N8�','g�6�"�2��wb��;�hX.z��2V�|H��������>�H�A�h��]$����cF!CL�0��G��,Ѝ��^`�Wel�w?�'N�	[f�s�0C�$�rK�� D@�|Z�i7�9��8�ϫH)�%��a����A"f���B�4r��"��Ldm�=��OT�zf�qĬ,c���}�"�ħ��~3�x�
A�,����Z�U9���.��b?��SH�E<�h���"\��8�%���.�i$#p�*�"��
�E�!�sz�ԣ��	�=���d1QO�W��#�uςl�S�=��Y<�.D2���ȰnO{a�t͖���o�-\b�    IEND�B`�PK   ��dXP��/�  ǽ  /   images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.png\�T����"  "%�R"��%�]�J7�ҝRҭtww�tI���<��]wݽ�Y.����;o<����U�GA�C���A��Q���u��y���s}X��y�($����������H����,{;)�z0�VP,~gN��,khm�l*S�6f��}D!3ܤ��VR�q{�Y\ÑV�]'A���fӵ4�ϓ��q�K����y���q�=~<I�����ӗ!hG{��%�M?�ă���w-&O���;z+8��Q���f���~O�&��D���?��e�yJ�@�-B�����z%1�����>&]���b��bp��W�	�H(a�o��d��-���Q�+4�R\�xWe���*.4�����oq�`��F8��c�L{p��ڢ��}
sR��z�S�!�����w�
^~&�*]��R�\H��sݐq�g�A�*�{��p���_���tcd�=㬖T[`��e�b�^Y0>Y��҆�R�L���y��up������$:�+􇇇�q2o��h�ۮ|�6 +ݐ����%T��0+�U����"���7��\��A����'��KF�R���������Jy ��a��υ�;�f��J;��	}|��j�b�i�]�|$1�\��s� i��~b�ͤ=,
�Ȁ��I>��[$�m��-"�c�V��g�~���'�����K��k>:,��.�"C����H��3�_$2^.<�U��)�	W����
ٟ?���*ȥI��+̕b����b�
�Tm&��J�](H��7{���w�xc��%"ҽ�Q�Ύ���<���Ͳ��kNtttfף%���qj�ES���.���8��a���A�Oԧ	�XH�?�����K���s� ȸ4w0��.��\�g�?��涉�Ȃ�E�L��/ڿ�q��1�w�0��ßj0�������@*����8�����E{gm�R���AY%ߣ���<,�QO}�o���04��=����_/��W��"BB�N�l��0�\@0~�h�U&H$�=��?�W��� u���YLAL$��Sh�,�٩�ha4b>�<P%oɁ�@����S����ez�R��M�/6��C�i.f�����oӳ�������S�ae*���r�|%�|%�MV��0"u�T����B�l���2w�$����u?I.�ꟆU�nn80�����00x��0�������CnbȚ	3y�6��7P�_,��
D*��{y��?�%���&PRVN�!��d-O��6�_d�����ѫD��,��V��c�݃�k˩�$^����96�
Ll_Q��z���)�����%��'.�7�ٓ����>�$g�_�1vm����
	B�^��z�t	
��;"$��UU����.���f�B�փ.��'�����뙓 �vHOW��3� ��S/
�����?vW7��KF<jF��Z�G��p�����V��GF�;�uu-7K�Ɉ�(!�a]�"���T�OM��<7�DE�待6���V�!�iJ�%9�f��f�����S�?2ޤ��CNS��m��^�?=�b��vjwZe����R>(���/�%�SF�'�g��a��渶�0n�C6�l���_����o���ͽX"%ُ�
����cka��,x�|t�|rE)Q���;��Ի�I��_[���W1Նp���eK�w5���b��k!0TW;O�/:"��M���{c�;�_�|E$��E���+�eE���K�k6��	+7�-��I�t�S
�^�r#^���Hw�k�����!��#�#�k�K%%�<\����D-���M�=	�F�dq�8�455[|�$��42�˖�p���c�٢Q��X^E��\�:��祺���Ĩ�sh��7n���sj���i(2T�E*aY���;�����LoD�Ă��G�����=S'owk���K-x_����>I�����D���Z���Ͽj9��!CO�7���{�K���dvu�o�W��aA�sbaqS)�1K�"�w�Q�ӳ���,}9*�΀���4[(���8��`��}�慀!.�?�XT==��0�*T6Ư�"�ڃΏ[���l%E�R'fH�p���E�� 4a������ײ�|�b1�c����aID��9wf��X��Ku�0���d�0��,^�c?_*��+l"�.�������k���Թ����ܽG
u.6%��M���
br��O$�N�?�?�bi���ܛ�\~�u1t`�0�AS=���~��3��e>z�����������uR�@�h�|Y�+�9�qM47��B���F8��&��O���\�p�}����uJ�y�H�k82z��_��9�"�5��`-��|&r�LS�Q��+%BŠrV,*����#om�.ל� W,�}9�@�p�H�����'����P�6�"z�6���?����aF#3��|8��?N�~{��;6��K���14��p��% ���8[r��N�Ȧ�B/��W)���e��ckm����"6I��ߺhwFDD�WEB��(qM$2)�X��E�/��$j?0T:9�TU��0�||��M��sC����(e����jZxU׷Q�
�}��i����D�۩a�� p��	�SvG�'<��ƾ�ãV����	MM︤е��Xp>��%G���*ӕo�"]�b���Õ�P��el�{Ԙ�� @2}�HI�X֦����ݱ11~7�;w�����YR���q�����&�����hn��,��Fg�؇V�S�^���>��.���4�榤}��������Ot�"+~j����"�%�`����W�
}m�?eT���u͝�_�Z&L�F��CDL�����9A*pkkˏq�pq�⡮���?�xW�I�v�SR�S:���J R�U��0�-�u�T��!c\�W@;Gj�p�Ic�tdd^��6��H?�v���_c����Q�C�� _��\mh�,,ts=��D=�T��_��+���_+��1��"�.5Vѩ�0�9�HW�
������NŰiL]��㝳��ԓ߆T�b-N4�X�!�ѥ�*7 N8h��׹��:���0�OOˤ�_EtَD�b��ţ|b'�
ޞ���QȐc�7�bq�b2_Ǡ1Nhc�1Kp�,�P�Ģ���o���F��� R��r�eU���mWa���Ƨ"�9��+k��uZ$�*6�Ud��Y�̪�a���W��b���K���t�<iק�)Y2�p����Z{[l���;=R�Kţ;|6��x�Â>��&�h��L]Q��ȒQ��W��\�E�����8>�A�����,`�E�� �y��7����YQ,�˧6&~qk/^���m�(�M�X��O������_�.s�E��L�n��PBv�l#����c��J�&�<������,������>ߧY%t���T�>�K������&t9
��چnA;���	����"����?]p+��hm!]��r�?_I@9u��g
G��\#��Z:O��0����5V?_|H��
v�x�&j�\ϥ�W~��s���z�ֻ�!����	Ve[�Su��梦���{����z��l���kr�V���s:����G�M,�<t����ю�a<`%
�g8�/�lG���'���n��.���y�y�0@�Ȇ|A��[���_cbR��"�pj�;�=iD��YN�Uv�����a|?<��1�+���ĥCA-�c�ig������D�DDV1�-���DMArѿ�_�m*���������²1X�M����X�t_����05��0~Ã��<��m�=;�M|�1y���ъ��݇fB���f�R%�Ye��4�i�S#�I�{�y��{���ȗw�#3U��~�#&���ԉ�ls�S�����Jb!v�Ϋڨd�{|��a��b<���0
��o���ajb������n��
K��gr8_f��/<��W|���V��20�"O5�T!6i[m��Yk|�Jhy���H!x�%�A1|*�v�C���h�h|j޿U>��Z���'��[��v+�bnv��@S����Q.J|<Mn�";�o��Y�|�[�o�h&ȩU��Tc�p,p�Z��ҼS9|�B�e�:=S�e�o^|�Or:;;v��I^��K�5^����.�͐�ު`�p����E>�á	E^�a���0~7�A}�e5�����.��\�dHu�3����ol��b����1tl��I��?��ҿc�ś�BQ�1(����"Y(��W�����=�z���7�Y��mN_5{�z�,
&�������9�\��і���-1$�ez�M�o���E��{�֎Kߞ��b��s$�J4�v�?=ɀ�N�:���Ԋh�J����Ս>N)�CJ�FW�%���iq�t�0/Z����0��X_b�ǂ��4����S��J(DG1ĭz��.-��ѧk�qpK(1Q����q�]X	�"�C��vf���*�Dy�`�����ǳ�!�-ň���C�/oq`��Ia��f�K��4�s�:�^7a:"���\�+{g���j�G�3z��A��+?������h��M(C��v��[�NP-&���{�e��O���q�!�9���>��>4�WX	*I7�;��݆���V�5��� H�*N��zB�I��}�Z��*�n�ӣ^fk��22�;�iqf���O�n�%����$B_&��W�������V>���o�Ҡb�W�&Xߙ6+I�RM(w�(A�`'}7���t+�sC;���x�������.S7R����eQ��f�&('�
�� J�&����FM
< ����U,|Θ�JM�_;�p;�;���N_�^T֩K�b�{AU��6�1�.5W|�����|��WX?��՗�|�N��y�lyk�V�����w���H�&��W����VS6C�+_F�}���5�ɪ>m'�Uźi��9X:(rJ)�����w?��Qu��!>T6�.�DsTr.jvt�|���k�C����\���r��~v����.�B�� �G�i�xJG��˗<3�vv�F�A�B賜a"Ga�_��ε4c��ɽ�:6�W�M�˵��B9�q������~=M�n��8�a���������[�P��
���uh�����A���g��vF��zk�/[��aM�������L�sR�ӏ�Rԯf�T0wE�3�Ԣ'�jl�;�0ˊ�=�6�3AuH��������0�7��F���XKX|E9#).'��FK��
װ}S���nǂ��,��jo`�Q��l+*�f�N��ox��x<U�����Y'��2�P��sɄ*��]SַHf�t_�!ى"B+ђ� t*� ����W������7p�_K�UU��Ⱦ;
�<MWZ�1�r�'���$��R�E����1D�C=�Yi1����U���_nC���	�d޲��?�h���:6�QJ8�vB`Y�CjP'8�̋���%�D<��2	������:V�`��<�#�<��P<uK!�$�Ԍ-��ѫ��@>@�v:��Z��n���a�̆ONl�_|��Ϭe�2��BX2Spn	z8H�P:��r��N@C/V;�R��9-S���|�W����*	�m���
��9���!�^<E��#9�%�!�qn�Ÿ6&�4zU]7K�yQ0��ͱ��?n}^�WW3O,�K���7&"�S�#�>�«���p6�LN���/�2Ďywtq���$x���S�������zh���@�ʾ��Ef�S�Wt��z�e�A䳴h��F��*���a�)(��
�
�mT&��M�o왧8������n�Aɍ8{M�6�Y[�u�Oq�ᵃ�A�׌�ڴ��RMK�-I��m���ϘõdT[��SW����t���*N�-�ҋϲ;��%	ג741[�y��h�"N�,�_P󣄗�V`:��hS�xQ����j�k9��3bCHԓ�{Oi��#{��dm�O��	N�<�m59զb��#"����ܵ�q�[g�x>�M66��ZC�h6��?]�K�X��c��ta�p4{Le1e�i3�<�~�8{���g�,
"H��Z-[��+*�3\��1���~/�s��K��Z�#qܢ��&�����~����,tO��
�0cبu/�(�U9��Y����Z8���һGBԭ�g�v`��$M 	/Ơ�2�K������N�ևr�ބ�1�ī�,�k6��g�^������c��%x�//EX�{!h��t����;
01��,P�<����.p/|� g�t��q�)���od��em_Y�'�3l?�熍���4�pm&cĘ!N��3G�ێ�����s�j�3�47���~�B`Ts�b,ω��-����s|l-��r���X�غ7:�G!#��n.y�8���)wSj��C�_�*{�1Jʟ��Nn83�sԼzы�ɕ��F��Z^���K��Q}�i�[  �l�$/m��D)�HH�YZ8�}��]~3�=�"
=@�q�����L2e��PF&�cr9q<ҋ��d���-T���O�����)Y��0a�g�ܟs}ρj��`�!&�mX~��u}s�"�M��n��#ꀺ*���}y������s��I�>%J���d�_#�=�a%oV5������>�P(�ph�˙?��K�rVm�/�Q�g�2?�e��gɏ
���xk��f�N~]�����hE��2*:XF))9#��p���bz�3�|�~Z����16���`uLL�_�����}��H��^���L�}��/�!Oo�?�Z���n�����kG�_qW�}�V|��y^]���t��Q֍A ��領>{I�P�c�&�"r��,�R�S�{�=^��?^��q��[fy?���k\���r�|��F�]�ߘ֤S�_z�6�h��5���S�v�qYzM��o�5��}k�noǙ���Y<�C�ƕ����/;�r�T���Զ������\9�9����}nH9^y�O{=à�'e G��|s�iɴ����M��f�_�X���a��m����r!.d��C£a�[x�Pռn���[�b<���L{���Oq�U�:��Lz��F�U�9�$�:�m��#��M���Q���޸Oدm��>n���[j��Q����k�f���6cbZ9�}CU�:�s�vpJ ������s���oƄ+=y���W�%Za��<Z��ڹ�/2Ƒ�K=�^�������gJ�V���A��v�����K�#�ߦP�Pf���p#U��.2�ϛ%n�TsNy�v��~ͯ�w��=�f[�p�<���>S�١s�|	I�&ˡ�P�	�[�\u$5��1߫�;5�������}��;�l� ���S�jGؙEzI���F��2M��s�7�9�/�d�BBr"bƞD�A�Tn�V� �}��t����s�)�
r���K���F�����H��hDov$ټ�,]l��>�9�+۠����z}�n�H�ȋ
��ʈ-j�"���qAl'��%gA0�ϸ���_���K�tt�_;K�*ѣ0�dh�2X�ęs�n#܉|/7�@ =
��
&��G�t^��:������Pa.&s�:F%!]�m;��pc�[G�'&�\�`���J�B�X[ִ�7ϲ�^�H��+}l��U���;\��rg�w2��[<�b�;jo���=ryCg�-���d;�q����)�|V-8hޥ�C�,�XVXH�zG��I�.k�4��{��Cw��IG�篫qK$�RT���oȴ��%X�u�2�BE�#!R���k�J\{@��p�	����(��j�9�|���G����Ifz���V�곾��ϒ:�Z5��n���V�܏]�ֵ�_�a�����lN�f+�d)�����(�o����C�;��Ȭ�0���k�	��_:&�lcH��ly��:�~Cn0�޶H
���\L ǁ���b( vlG-�w��,�������_�<�����m2�;���}�#C�v?���9�K;6od�mH"ÅV_	[��A�|��l��'iD|&mn>S��j޺�����A@��M-ox��v2��߭0���v	���� Z�՜7�dnP�7�|r\
e���f�F���I�>�Ev"Z�$�e��9�O�8^[c@0��0�UU�l򎸟�"����������酕ge�/�Xj�q�N����X=;#�����rP9s��=
��~F�U���q�dd��Ё��o�����v����ԠayRjU�[X,Q�D@�O�Bd�=��l�fF��u#�� 6O)��%���_c+4�-�E>qڋm�������8� <Hd�߼ϕ�Q."q� P�s�pG�	�#̇�wq�x,�Oi0Ϻ��7Bf|ۺ����*Z��+�eQU�";[�=���f;�3���-< �E���p����( Ԋ�E��J�]����ec]�B&�++6D�d@n�p�ĄH�V/����9`m��˕�F������hkk�벽@���<�
ݢ���aT�0.a~���V�"����E��iPnp	�ǭ��beU��+���ddH/��I���?K��N⯢I����DU�eR,*���8(�H�j�

&���~�c���՜��7s-^,3[��6[s7�h�,h�5J�9��
���k�*N�����3�P��)��C��`�nYD������w�CZG��jk3�j�������{Wb�4��`I����B�Vz��i�����5����G�D�t1J���$�f�5w���M|v08:|�����t�7��p�A�R'�h�d�B���(AG	����-��-\�FA�b��j@BԵ	
4�˝�V"x`kB��]��>)��;A���0��A߶DZ��t�@C@i�C�_�*��mmS離��i*��-���qI��NS��Qx�����>�TIB4EC%q
��=r]>&j��Oh<�u)c3V�lb5�S4#:~Q���}�F%���R��u�DQfG�Ǻ�B�<�c��	�1��^|�r�v�X��w�3*��V�����BPN��<fY��=d���U���S�1��t�K��� �Q�l��J����h-%�CWH�~!�*n��v̞��ݶ���MP�ٓ���h�i��]�����Mg�ITÈ1#XX|v���j��lE�r���,L�Y����6���v�g�������D��bK���J\�M3���q�H�~a��Rx߾$�3Z��Pm�slӂ�O x��G#����u���A�L�����F �C 0�*����� �]�.ߋ���E�E�:]e���R���y{�2��Όߓ��x._�z�At�f�|������'��!��/�%4<����-S��A%��冽y�R@�d�rL��5��E��BlR`	�|��5R�^�7��l�1�w)Ӡb}�0���GD�}ng �Ɣnӧi�F�l��H<��j�R d��$R0�?)t�1�=O���7^�╍�2k"��џ<�L�ݿ�Mk.o\�Y[.��jY*������a�M�M2ׅ�$�~!�	���0�Gy����]�br%/�|��^;��(�� &^�<��1��p����Z4�`��F6�T7�k��G#��p"�D QFz��j[�z7�G��n�cpS\� ����&^� ���aM��k�D��v*V�@�mù�("	k���BS���od���q_?��9획����OP�B�I��+rY�(�l�:�����zL�"O3�*����qZ|��u�/f=��`�b��@æ� #q�]k�?a�)~�򶱄�h0j՝gǮ�#vIdShIs,���˗����A�PDz$�~�%�����p�-�C��G�����w~Hbn"+G"$�w���_k ��[d˻�����a`l�����_!�����Gf~0�/g��[���	AT(�jú�(�U�l��g4��ul���+��^y]֑ex5��nLpǐ \"�.���u�RYLA�, T�3.݆��Z�q5(F>(���:�|@��ٵ��}��[���LN���
�g���	hh�ҳ��t(�T�HI�)9Wq�����ק��IP����V��ܡ!!���!:,�1�	�B�zj6�^ ��c���I4��x��$�4���O�k��JG���@ރ���>�K���ӈʅ��B;u��{
/����S2���B/���{��	_n���}�����
�d�T��ٳ��?4�@a���]��*�(������O���T�ȑ��`�HU\=yr��Z�X��an��CdD΂�����4��5�#J�5C����D�48I�]r�n��r�x,�
u �4�w4x��"�X��S��*m4W8- ��$��+����}^�.}���"��l��S�M��pP�N���H��+�B�VbKq��������Ҕ������n�.��R�b��V2@G��=~�a �\-�BA���b0��>��� 1���5����A�����sC1��� �D�;�7_ r?m�4��~����7H}fx
���~��Z���~M��9��.�*�nk�x �5;�&�y��*����+�`�T����K.��oD��x�7$�ut`==á�b��R����t6P��Ǐ�B����q��]��'_k�R^����1Mz��z��Qf)��E"����4��C0C�>�<��yE!���rK`Y*�=�$^����T6�Xɗ;�%�JA[Ԩ�[mH�m��Ph"�-�$ݗ<�pt�)H=)=:�d𨎿N
1��߯ 0�Ej��\�팷q�q����s��p��.�~�b�y`Aa[4�J������"Te�CP�����"�9~���=��g��9Y��B��[&��Π����e�o�����-�3���ǳǾ�h�UE���9�
�ʐis�Z)�#�-h�W�� '��]2D���&���Gƪ %�02sr$��(i�d\�
�1ެ5����(���X���ڟ$���T�li���X
�R ��"�o�l�FrPQ��m>\�MW����l�cn��e6YT����_I��8�����ⴊ�:���)t�tj��"2�J�ۗ�ǃ���������Hl�K+~@΃�Wh}�Wa�<�4 ۿ�ݲ�3i�"�C'*�DT�^i.ܱvۯ���>�0�B ���z����=��:C嗣&�&>��C$iy��>�<#;x�vwե����@�]x��#���<孷���j�x������f� zX�S�aB�&u �z�!�V*�$ UO��b�X�Vf/�l���%�alBF����騜U��gi���>4�kjj��Q~92�ߒ���HT2�e�.�X����# J�s��y�l@�4�. ��4k�&��>hd:� ��6H��e����h&��c�T��b�9��t;#{���#��y^J$n�h���z����J�uȍ_ݠL[k5�e��qH&zn/����A�|�����������<��a>�ջ�l�f�}��py�.l���R���j����_8XW>!?��$��i����s�)Զ�u�+o����6 N	�s���ɀNl����l�jP�K3��Zt�TPnj��g��9G덊@e�(x��[2-�HY�9�Q:�I瘠��:1ǫ]�G��0T1�T�z+��zf�鿻�4��٫8��K�~`�F
F/�0!"g��D�����}�5��Kr���3X��	�2��uv�趆��S9��A��Q��Ȅb�L'l�d���~�]Ҽ�t3�~��O���.�>H���>9�Z�j���l���c��l���؛zq3�O����f��o�cي(+�~��gVB��2�K�)\d~�HHA���|�T�%^
0g`G�Ĵ�C,��B����[d��e��w����w��7���1mh�2��f(���Y��m��xs$����9�lr2��-��!f�!7 l��I����N
D�ٽl�7�K�Φ������oV��� �<�.�*@0�{��i�E�����\K�meߗJ����]��.	������?RPHHIHII�ʯu=D�XMՇ��ݑ���A;a��!�ZG����%Wi*�;/l_֐R԰7 *$OE1O�A� 3�&@M�
{�G4sds�]�a�VE���
������l��� �>�Oh��eyPJ]��]��Q[]�,��o��b��v��<:e�-W�Fɚ]��[�a�Ҹ9[� ֪�=��Oz4#�l�lRX0�K�1� ��z,�4ğr� h�V��� ۏ�"�-��v7)�Y��zRH>`+~�wfO��A��#*_|�7��wbc�I%�"�h^`5Qv�{�б�����8�e}����׸#h�/:����t냆�ҲI(p���k'�&�^-���H��<��}o'��S�t˟tuu-I�ɽ�ɋ�P��@��v<C�b���8�j��d���ː���w�j�4��ٿ�L�I���m0$;W/�1�@
A�V�p>2<,��H+<-�Gl��hM�'�f�)��b��N���#4m���8����B|���K&��t�8�"� 9�L}� =�i����+�b4���\*߫�]̙;������h�ɐic� f���\H���0~#���:��[Da�9�hSq(�Ua1��R����1����M}��@�5g�&� ��m���'<���rn���oR�#��6RZ�룠9�!Sex�p�C�[hwh��UX85'&���'?�����$���:x��vҐ݆�mG��o�H�|E���"��X��~��l�``�@S�����h�X��΀K�$Z��s�X@���U�H��br�����E0/!H �`h�3���a�ێ��O�j(�P��%6O��IE����J�� �0�p�n��u&�Ā���*�}
H��_ł+!�m��݀��*�c�@�+�7�����l��X6˭<�;M��$�n;�e�x�Z��g���ԧ��Il�+�F�m]rh�� 4C@AF����a��6~8
�#`f@�7�)\0���4���<�P �$��X狈^��a��� ;��n�"�l���-�yy��G�dn��� �-)�~�r�x� ^��?ˬ�a�i ��Ѐ���L�138����4�����j�Ρy�l�h^��������	�J��6��Hb��!���`F��i����W�7E(��Rm>��� ���^d9�p(wt䙙~�LGճ�d���	A��ܮ�꽏�����{�;mp�6l�R�1���2��_{e�Jv���(���{ ,�U���!����)�X!��ܚ�(;�~�2!
�����Iyq�E��ݍX�A���C�sw��\T�d����~���9����5�)�l`��90����כMX��[���r����"�#ض̆��r{:����^��z8��Z]�r>��|�
���J��z���ɝ�H���������_�X�x�p���>V�3q�S�WP�T��S�����v����L��f���wu.��V�{�v� a��������g�L���gVi{��,�X����9]K1v�����κ��l,���:��.ju��d��&�Ϟ,2���]!���i�.R�U�i�B;�mFf`�+񽮸ѝ�u��q���Fh�c1N�n�Ϲ|;?���b�i�n}�	���,c����<��O�$��|�5�ި:86. K��I\Q6�yc	��o�r�(hIƅ��A���W�����}}�㥠=.���������m�M�
?���;?^��U�G�~QR�����Ix��	�[���+�_c���8!p�9����y_����cp�j}��p�PU��if������4}�������y\-X~���Q���@�ɝ���+���_j-���#�.R�о�[mkݶ���P����G߉cU�dBǎ�����t~*�_ʨ����o9��M�� �g��r�w���5S�xd�M�����C�zǫ�A��k[��w�H�Fļ�h�Iv2�^�U�+�Ľ����^��00���k�׉)z�F�UI��F�=Ӷ�׍hw�=���\��5dw�v����Q,���r�����;)���� ���2���i[�E{�|;�5^�����9�)�U�-��}&ZS��k�z��樿U^�~�dp�d�r4��u{CJĞ���v��nG����K�����:���@�s�{G7�:���v����ކTW[+�����Qu�[t�I�jG�s>�X�ٮ��8�hEn�~�pGl}Y�_�T<�{�~��\{Y�N�&{�� ����dx���Hq|��w�_�mџW�OZ��%�=y/%�;����W]t:���ӕR�ΰL|�'��P���r#�-F����5u��7Ew{A����˖�� ��yΆ蔲�k�b��}�xû�����Ҏ)��\s�q������ֻ�ޮ}7������:��'Qt�V�7�9WB�O��W��s�.��Km4j����lfD=�MR�6j_��16�-���[�v��7�ٵ&>1U.{��T��AY��u��ߛ�%�h3j+�������'%2��:��X����kk�����KB�2�}s�f���������'k셣k�4q?�8���J�l�%����*4���6��aN���6�P��<wĮ�� *����*7`��$,u~�p�&��=���B��/�;"}򑢵����*=�{�|ԅg#�Ѱ��-���%�$�H<ߓ9!�fd߳.ץ�Y�fd�W�$s{J��AM&	pG>>4W��p��k�DG�l"nsE�8����f�M���3È�' ::����!�zafn!p U.�������f
�=, �+y�e*zW�g zqc4`!O�Gs{��67G����z�&-��r^J���+�$ex݃� 6�_��;�|�}|��wW5p���?�;��+\Q�h��K��L�N�|��滸�5��`!�޾ߴ���d����l�8�V�{����W,�]]��u�����(*	Z�o��NQ�9�/�g��6S�ÌA ;�fM��3$`W��\=XhQ1B��m{�=�:���$z_\i�{k�E-�N�ɣ�����,��:������L����*��E��;׾Q	�� ��(�8(�G<RXI-�S��ߒ�6����4�\��j��|����CL%1�,i��J�sP7	����>�i���R��K����ۻ�M�)�g��p�ܟ$����~�/���z�Fݥ��HV�Cj1@
�]d����V�W�I��l�X�
)�np��\�l�˩��oT�aaV�����	9���Ȣ�~����`9�Ǧ#�M�Ǯ��.BYu����������cH^ �74�g ��eEFwzb��7\R������W �$-��κ�D L���%b��	5���n�&�[Z;)�$1 	��3A".�[?��
s�^;��/�Y�@x�VR�����0;��/CO����1R��
�Sw��8|U?�b��g�O�-!n�p����灒£�?����5��fx��4y�g�Z~��yU��`n���=��x�>��¦�*5M_6�﷿�o�uO8u��OuE5樜>b�94���+�n8c���+R{��|�V~N��j	9~�on��ڃ���ѝ��Jg��(�%����]U��yGc�[9`s^nJ���'	Ԝ��6�t8�Z�ޓN{��6����,*~
�̸�zƛ���P�H.`Dt�vBD��^��DI���S���-O��PVڽ`k���Y��C��Ư#��w��ʮ�u�,�P�jGy��ߏ}��ke�O~�捎�6�5�)�֢����zG���֚�����B�r�"XQ�o��uɅ1fXo��PX]�[��7l��pY��6�I��w�i�z������v��J�%婻oa�E�=]�.�~�G�r�?zJ��4r�H���i�00N���#�,Q#·^n2����6���8 �$B�@�L�}�b�^W��(��}~��dZ���s��Ni"��Od��I����%�8���/O��/糿���?�sK�~w/a�e6��U.�"
���n�ϒ�hh�b�a??�\���h�Q,zG�S��`j���)�~��
Z�y��fѺ+����#ꆸ5�ݤ"������sLWy�������qP'3�T�F䥝����(�4��X�~��l���ğ��t�,�V������]�����W��G�85M�.�F⟠�heU��p��}WUK�?�ե������P�U_[ˌ�v���.b�+n)�n��<�]��?I��$�@�V����uճ�(�?~7��L��uX<�p��7�N3k15Wk�[��Ѿ�k��j}��Z;n�h�?�н��8�e#���+*ԏ���Y��/��N,ե��ȼՈKm�G2KҎ��������3Α��?��SRo x�j&��Y�������1�����\9I������Z����:LPЂ���"�>U���	�*�����O���'�ӛe�y��}�Km���gEX<H�w<n�8c4�eE�H��������M���XZ^�֖���=�3��P�� |��������NI����ZoT�G]��kn�6�t�ܑ�Y�����g7=��^!�늀T��Oq�s�B����$��l��c���/����,R���ѼՓ�]����>��3��(�[a��@܎�/����N	�3�}� -^�h�x~�� �Q	��X�%�/)�D���ao��S����o�y+`p����8��Z�΄]�ُ�؀�:�%���6�.@S7��G��H��.Ȍ���<@�J��e�A�>h�#�'�7�;�ǫ~�<���+Ϭ
_\W�~ݬ����'�~ʓ���l� @dx�uk莑�9=�]�v=sH�����m�ĺ�%�\����4w�Oy����g]xz��48��`�[�nI9��z
,��׮�]{�h��l����o���v�����޿�~�ޘ>�^�Mx��i����W%��ȍ~����p��)���%Ĩda�'rh10-M:6i�� cfA�)%5���>� �y _/ ބ��N�o�1�r�dg�o�|V��5"�ܗ��]�k$y�2Y�Ji>�#��A�.6�H���_�]ND�H�~&����@���@X�����T���c6��fܴ�R����\�)�C�l����z�=��QT�\��V_�x�죵����i�\��.�,�f�ڽ���2��"0����&�Um����T�OdL�S��dmMU�Q19��(�c Y�<����<��p��w;��C������bzV����|6z��Z�0H�AW!E,�8O��Q�F����Qƪ�&,P9��9ƠkA5���rG���W�f�r��y�jp*��~�%��CLP��A����|w�����^��+d�C�~�	?%��d���+e�2�I�����o'VL�U�M��W�?��d�]�{�1K�i��J�~8��sᚳ��s����N����h��{�ㇵ�������{�QA%DDZAJ��K��E��`�!DA��`讁�������{b�O�/��Ď{_�u_�ޏ�E�WD��Rx#v�n~�w�I��)��tR�m�}��xFj�tߴz���,�%.�[�@1>�.4~�-��]�g�uY�d��؁���|BYfB��?�,G��{Kf��d��IG6���(g}����"Sީ�t��eyGz��]]�^�~.[AAM�I)g��@k@zԥD�MQ��L��b���c�D�`_w6�U�f�����9�޹�ܪuW�}���4S�"�L#��J�#!Y���r��;>O:���E�%=��i.k���=m�@�1�ː��:46T�@sQNoma�^�M֔��i=�a,��;h�AY�8��M��@��pM�������C@R�j�>qZ�j�$�i�����<h���1x��L�pM�/���?��K�(�^^��T��r~18��~� ��#�HƵm+��F�: #ؑ��0Q�6�P��)���W)&l�_MT��,�0!`kG��^�������w�����i:��,Y�]���D�(�m���I1f�K���|!��"�e��ȝ�	'�WǵU
�r�ɶCЧ�z����@2d�3���BuV�n�}.����]�1T���8Ʃ&k�>���Ī0I���ًY�l���9���wQ�K˔=��-�x[0�6��#w�����KX���_T�f�S���i��#����_�x���(������O�~e���<������7!S�xSd���B]���B�l;/[A�;oWۨ�t��ݢ�����[ߚ7���9>��24$���G��O=��D"�Yyޛ�2kui��b�׶c��?��Iې��yr&��&uT</ ��"�o����7�}.'�j_W;��H�1ez�E�)fd�E��	�͋�)~@'�ǫ���z�Nļ�!j<��"�@�����۩Ǜ�i<[��_�}�J渗��-+��g�"�Q�vIVWF������C����a����W̢�Z�|�&#�p���X���rb�˚�=Å���e�	��'�Q,L;�[�2�_uE>,����}�=�Lg
6yx$��4�$�5k�A�8�|���]����&�,]�c�u�w>����.�~�ъzM��bi¹[��R���d|×'��(ݽ=��䡯�b�����7N�)~�I�$_<�rW�u��划ĸ8��Tt/w%^��N���A��bs�?}�"�	x`�ř ȍ�W�����&yDh�_��:n�����?����2�`��Rx���-G�S�Ǩ�L@�Ȅ��i���p���S��@��j��Fz���Ț�r�P��;��|�w6ў�r�NxkBN<�Z�NtP���$�jvH>�����~���`<!���ne���ځ����@�����]�:!B�1����!�s�m�Y���r���È���mZ�Z_�p}t�ޛ�f���9��"�Ғ\:�$O��pg�>v����k9/��B���E�k��Ne ��(�`v�E�$wt��f^�]=U�Ć�Q�S��g��F�ٳ�y0��ލ���h��1n�
��N��(E���<��7~$����b���g_O/f�N]q�hH[���M̆�# ���� Ͽ���]��>/���%����EAF_����)e&wa]hI|h��eߛ���gKk�J�mׅ'������ќ�%�PO1��g�@��2�J<m?��F�7��t��I0���kLdr�~U)`s�E� Ѩ�{���jIɉ=edXʓ��.��jq�����Ͽ���xH4�ڨ�1��p�V7FO%\�!�E�̑�1r�3`4/h2��������Um��)�R���ߢM�_�}�S��Ҿ��kbN��[�T�>�-/z����ђ'j��x�Axη_��Ʋ��a�a���^V㔳f$�h`��׍�����q%��jT�L�J[d�t|���*�z6'�db�/(�'���d�d���7�`:q�e�R7޽[�ʲ����Ҧ'��N��#m5"9���0���ߠ�\��KzG���G�Q���F��b��Bun��Rq�J��s1'��3z�(8b2���R�`oX��q��
ὴ�k��Ϳ��?o�a��\�3ct�a��Ez�/�P�(4���5�S�7������]�>�V�T�+�Da*腡��̊=N(��&��8<H���Mdޅk)�n�l|{�������{~�����[���y�X>Y%�����Ԉܯ)�I�\'I<�Cwv♩��BN�����b�ĥ�]A��#Rb�6���[0��n^�
��r���@�)tnӛg?�H�{{��I��/ͺ�`T~�ۖ
\ڮ�-W�|r��,핿c�X�哗~!���nS���ܼ+ho6da^���4�#��n~O����K#���`4%��溧�8�Tm��A7փ*�5yFV
[����Y	i�ya>�ˏ�4]A�������Hp��i0�YE�{��,4�ڗHf����LÈ��;,�� �J}+OQn>�gh��xL��X=���{j�+#��ry�]gՎ�rO���f��BF�|Ԍ4��H�li�e���%�;7�cr*��疝I�W�or&�8A���+Ku$;��7�RO�ao��lr�!	�|�d5�몮]y�ѫ��d�C.���;N�'w��l&�v_��{�K��f�S���/����WI��X�r?!=dM���X�i�.�����I^�.Hg�X�9��rY�+�S��T��g��L�wc��EX�MRV:������lr,�.��M���3N��W��t���T劷�/߾Q`
"�%%��S�u|���{b+���/�dz�6ș����ʓ�
�e�T4�J60ٶ�$0F�#Ll�C�\��^a�,1�'tҖ���Reu��mn��mޟz�M��od�7)�klu�~��_�X��4/�������p�D��u\_z���I�W��DX��HWl��rto�o~e�)�lh�96�$?��F�^@����م8/;�ћ��\�k��r�<�m\f�y���'C�*5;�:��7I)����
qtY^�v�X���<�� 'B�1�V��w�{s�e+�x��+��TK֣�v�e��r,<=�$$$�#�C3W��m����^�����J��UD&}��������Ok񬎑����+�!�dU��Zbo3��������U�Ӡ.�@Tп���?��n�������?Y�n�w�i	��pI�q*uv�*��	�l
M.z�"U,l��c�l�}d���6	Q�#QHv6q��.��Y�daN/]%\�k�F���[��:�$�K�����Fn��Yh�b�F&���.�"޽,q��#DOm7�k)���6��Q+�L�(#��(�Hg\y��VE�H�S��'�?ޫ{Sȁ�I�S�F�n/N
��&�Cf�ɷr�]��a�_,U"�^��Z=��r>�<+z%xr�X�5�0&Ȳ�����p_`��.(��o���
���â?��2D������7�V�/�����_�ܸ)o3k�n0�>���W�8�qB�Ιd� ۆz
��	���[o�T�UK�o,��ׇ�v�������W�,eb���W
9X��%�b�aϞ^�"�(�!/}�c��&��M�7.��|n5�?�F-�E;�b\_�*�蚳�5.���p�=�2ȎR�ݝ������z� zk1-�y?�+�E��a}
EC�M�'�n�+^��3����h��hA��ُ���>6#[UR6�9J��D)�19�<&�kC�� ��ti~m�u
��X>�]:�mۏ*��_$6S�9��?���=�k��N�+~���o���*�53W�ޫ8v��L�P�с@,�����h��jج����
`dq��8:�s;�=D/$的<�*�����JTW�y�V�* �-��1�H��29��M��(@;���� ��4]���7��w;v�,	�9��}��p�*<���p���˛K���89�����u���7��I'_Zjn����ʖ��������$+{h����tBI|Lx�ى�r�W���˔�P��$?!]=���MY�F:泰�2�>� ��Du�M�tb�rr�VnKW��S���,ƕlUفD�GS�;۸�&���������5�5�h[H�^Q���O�fMO�-J-(J�ƽ��P@ (p����ξu�V��~5c��/�ˬ���f����v�*w�ᬩS��=���}���?Y�q	��U֗Wg45�P%�Z����]�p?�����Z�~	���i�y#����(�~�y��K��^ڮ,HB��H�9�|?滹���s~W=�m�$����i��Q�]^5z�c��V�'���r�p�^v�5�z������>��)��|��(o'�wR{�o��8��IИ��I�r���ξG����u��ۼ�4�l�0�+��	��eD��=@���V#8w_��?*��_���7��ųr��0�������>�Ye��WTo��x��1��%�� �(�`�z��/sI�D�o�V`U��3N��쌉�u���5���ŹĄ�?�BJ��~���ؕњ�;2��Ns<�Z�y�i���r�_�)r�~��n2�2�SC6�$җ�b�����t������(�ו��0(y�k����덶Z�H�
��'�K~(!��]��-�h�(�I|<�㓟��H�$���{y��j�����-CȄp���[���Ȃ��"�>����SX�\�����N*Q�ȴ����b���[؞�����]c;��I@O�����0�̭�K���Z��&rٍ|�JXc�L���-�<��t���L��������8Zۤ0�y�~��"�Ef�ۼ�xc��r��<�̬�ץ���q-�(��\nc���d��I͟z�4 �8C��篸tH��/�AP>�ii��0�I�SWEw�������j���(	M|��+���})Mr�\\�\q�}��ȝ���d:�{h�V�.�h�cx�#\��b#����|�+zCB�[+Ȼ�>���W�G�u�LT��)��_A��@�|es�n/�cut�:'|���Ǎɺ8�~@���zP�j��ρ����׼�O�b�R�c�����Y����	�o%<{�|&Mwo�B��|�g.d���(6 �9��i�!h;e��KbM�������"�ک>-?����t���Y-�=QQ�4����iN��7�(b P�s��ݺ�����fe٪��h����H��Q��ǎo5�6��^�&�)�� �e*��.���6��OҨ]���0��#b\� �1���*�?̂�1�oS��ϫ�?RB:�.�k��yR��[�s����=��7ys��rj�L<풐6u����zn�>)�SlQ���_�[:����uq����������_�,���eH�TB���.!|3~�������e�SB<h�`?��*X�7��3xD~;{�<�M��M�0�4����/ �qdޟ�ؕ��W:�'��ZIAϙ���hh�����2�"?n/�!#�������Ȅ���>�ގ =�- X�է#u��_EJ���c^�r��wA�	�$ê�>��J2�.)��L������`����l8].�֪��[���7��W�����k!1��v�u���X�=�{_'�X�뷓-C��N����g��
�U6?!�Z��3x�&)��^'�����xFv :�/E]��_k�\�������S��>�9aF`2�Q&i���_�-�o��mR1KS�5Сٝ�	�|����lO����r��Xu���>j;}�����G���tBE��	�hzP�7�@�i����]I�]K��F��̭9�W7��]��3h����}��mKww����SE���Q�w�/ۉqv�\K�b8��è�52��=� �|������Ƹn�w/���hD���	��x	}w$��MG�vko�Ę2m��7L�t���ӿ�Lս;�t�RK�&Å�t	�I_�ʹ�V�i
��������V��x�x�jR�f!��~��C���̇�q��0'�������a+ϳ��})p/���U@
ܽ���<�
b{ �V��-ZB'Y!�w8�v���A"�p�T� �D�w5�+D��g�[��۽�Phཅ`u�Ut���T�'ٯ���- $�K�7)���8B?HĦTﺎ+�
����7��Ueܭ�?$���p���~��r[�W7+m����`�ω���@��4��;�ܚ��8�1�ʅ"��v��^.�/1YAA:�6��|:���

�~������Ns�S��gϺ#`"%�/�� E��r"�v&^��?~�c�_8��,�J�>%��.�q�����Ϝ��]�� Y�-7��^���Zz.WZzl	��ȱ�\�b��è�uC���s&�6�� ��=|�R������@���
r0�lu��IF�?=fb�R�� � WzH��JV:7�E��q�W�&�Rv"v;��;�3����Y^��<�.��(��@�䂇�F]�J����f�?@w��(N���k��2r�_�� +��,�С.�q~о~���V���fN�6�����NG�'ci����VR-`㸫���te�Wg"upɣ��Ke7�ؽ�q"W�,p����ʽ����b}�k�H� ��C����\�����wo�Qf+4��"�-���K;5��tq���c�J�|�l�Q���Y����t*I-H���zO�l+K��h�UB�c���ճg���\<�r�rS��}�H��n	n�U��~����b.g.��je�B�F2b�?��%�n�\�tV��UZ�@tP�Rr�ټ�!1 !b&r���Aů�>;�ܘO=�'�_<��p1�������ݐ!;ܪ�vn��80h�q�m7�����>��!lW��kUk�<̣�b,/v���`��S[�:G+��P���F'w��c <Z.X�f6�`1!wْ��Td�;��O۠}Wp�EC�~U��ݲ��UE��z��7��/�?M�M��El���C����e�� �� �|8��!f\��ʇ�J��aѷ+?����M� ���1U��EXCsপ�����;�e�Q&)}��m>�w>2�q�����C_�P-�5Ir�]�o�I��[�!���!y�ڵ=_iқÛ��w�Ol�VI\��[���&��C]Z�;��=������^С,�à*A��>`�?
����Ʈֱo��^�+�.D]L��ȔM��C�*@���G+�즶�ǒ_�.�O��{}���u)������Y{��(j�c?���u���c�����S1���^���W�ٞC�ղJ"^�6����[�����J�2��z)}`�j�y`a��4!�ck�6�b�]�x�"+{-A��zNr�"�\`2�}u����Z���t�\��k����i������2\����֏.��	�����r���������|��}�b��8xl}��u�
YNԪ��_B7�(<�-��;�^Oc��^�������O!��<uD�C������8��hB�``�R?�Ҭ(@���q�}MHh}�W�δ/띜o�u�U�+I#�� ��>rR#'��#G?q��<G���Kt�ޖգ��8U�����&��^.�C7����H�PT�*����7m�M��X�a��x{�����w��o�IFHl��t;���qd�]
C>-Rg�.ebe;��D�o+N-/OE�m����m�Ȃg''�3��v,��0Q�U%��6���c(lb)�5�ϬXBF	�.Wk��C�!���*A�j��č|P�]=-���^+:�NK�T�#�]�'���q{�d�L� ���VN �����>=��*pc���Dw�o��	��0o#�X��<j��(�A��B����U$0C9F'���ǝ���u�jO�N/���rYyNɑ-\����Z�d
;��V�6^דv������=!�ǝUȔRW._{��t�C�ֵ�/�z����#������Z���{�.���<M��*|��K|Z�ՊƝzI�B�<k`I`���wU�7Cu#3�%P~��@�XZ8"�M&��f:v���7�Τ�;m�������!�u������]2G�I�g���+���E�+j��t$��{*���=ۮ^����@ł`��Y��,�s�@���}�B�� .���������v�nB��5X��Ωg�9��*Gi�{�9fd�zt0[��x�`���ê������ȫ[�X����-�Rv$�Θ
�����_�H0� Y�r�_���X�D��ݻ�Ϟ���(k��Ctө��.�)V��3q�uEʢ�f��y����K�+>����]���SQaR��KQ�t�ʇˍfe)�T}u�]�r���`l�ٕ�����Ӿ��^��ʗ~���㮝a���c��z�xX�,_n�[���ss������A*]���8�x�m����7V�ը���?].�3GBbJ&'��
�MQo�Hh���8�}-�b�n�O3�ʙ
�4�>�G�̀m��g
�.��H�):=)5�c�$L�����j�tS�f�R!P���#w9U��zNlU�V��&�ʖ�/ŧN49�����E��+��;R���nE9f�����H������:�"�5�1M�x��Ѣ�6N�Pf��ߚ0�V\����p;���"ʀz���m�1����_���Y�MY-��{d�H���x2�v�n�m�4�X��s�������-W��n���9e��|�������.T�k�;�O,�[������o��k��z:�?{�m��YXR���<��K�x]�e��eɛ��s��r�u,:̮��)�'#�E��^��J�aųgTd �`�^ǻ���Z����D�y�`��sz�ۣ���g���`�V�"��Gz��ꍼ��̃
a�!����AV�Do�-�j���RPǱ��}���5ŴiJ8X�5t
E��&��t����]�R J&��eka���.���.e,r��X�2RօҴ� �E1)%�+*{�����:��0F��%r2��-	з9�7`��A���6^���f�-��p�$x���:�*�w>Yb��b��"�4J!��30{���L$GTF7\�e�JE��z}g�A,�O��L�f&Vd��s7���/����c�Ў�Ȇ0R���:�2P�y�����7�Z�&�j����
��������i��S�`_%I
xRC����hb�l����~^~N(!�\�|��ߡ1��×��A�^H�>
Q�?
�5ղ�Y����/ 3|�8�
MQj
�?�wS1Ў6��Nme�G�҅]=+�r�.}�d�CE�bQ��������0���/��S�o�񥚡�1R����?cP\"��79Tc���b)�M�k���ٳ#g`�q5�8D{�(��S���Gps(kDF��]U��C6�9�+�&+�ψ�s�k��c��0G`r�U�=D�ִD�^�n'��-\"��?5��>\��0_��N���U�ږ�ls���E��+�K�~/��Ŗ.��O!Ҟ؎snc��K/�]� ώ쿾L ��p>�Y7]�����#�q�f��O��	Ӓ�hJz�e� fW`��*�� ��,����ʟ�D_
^# ����Q�_�m�/�v]�����X�82�Q��~�f�2W�'��^@����������ޜ{u`�:.��i�z6��L��
�w�,��U��!*'��%,����]�\�{>ԋ|w�}�Bޟ�=���9. �ݝ�-Slo�+�3�^V�9B,x���x����d���5z_-K{��lt�	#J#O�ٗ�����e�~4��v9�,B�:k�IW�6����r��k�voل�*A[B^�b��R��v��e�o.����N�QV�B�,T��LF�+��u7S�QU�BnS��ߏ���nɅ4{۔
�=Tƭ+�~u*')�W���ͻ�?�m׉kb��`���+j�yŬ=���r�[���3,/y�+q����F=���T��J���3#!v��(K�m $��If�8���L�E�([J����[+S�����
��8f��޾|��-���_����a�ź�({:�(q��D��h7?)��ЬtR�9��V/�%vcZ8p���Jf�r�O�D��q���m���3���)��;�_��P�U�`鵰�u��n��l�����7�����zUTR�%�?kB&#�gݷ� $;����xX+W�ʗ�AO��//���Xߕ���p���'A��]M�	���~���q���z+���{#^��h�ī�g�����Ɂ;͗�%�� �"*�.S.kXki���Z�1��*w���-ъ鬌��P7��"�U�,p;����h�<-%
j�].4h�<�Qh��- ��SN�T0��Ȥ2csOӴ��V��_�E�z��6S�SH%�>�&�� ^h�ѻOx���ֹ�|�&O����M�`���Ų�Y���߯�w��C�}�be�w�yz�E��"atP!`L��P���Oυ=���~������c���@���R���o�Y	������r���X#�6w/n���D��pL�v��f�8n��I+�fh���9�㉦�鋯�x3we�/���~��\kR�@�<��$�|���g_�+h�ˢֆ���9�g�?�IXQ�R��������1�%������!*�t��_޴�L��}�(�l��'%X���;sBx#�ޝ�^豬�'3��T��/(\���P�K~T-��Y���y������[�X�
��]��߸إk�g�V%�����S��^1X%��W�}��<��M�"B�p�1�s���i�x�h���O0}�c1��{���b���@��Ǳ���6���E\`0d�\)mqF��#�f�������4�����ZǲИX {j��p�@���ecY*덾\�}��<�T����g���[����9aa�y\J��U���(�v�W/k�,lx0�.?�%��|Ų���gMZq����e���0�$$��2e�8"�;"�,+�-�P
������a}{��C8%nr?Z���� JKN�S}h���p0S�������������{�)B�^����HEр�ۗ*f��u_�V}@��x識	�� E3n(����Y|����nj��!l�Q1/Z�z�4~+�|l���4˓��n�qKe�(� �Vd��;��S_���iM�"���v{��=ܬx�:b�g���by�I.�X�n"_��Y��)��?�`�Ih8ǼN�?�#l��i+]�,�,�~�9=���)���b�w����N�?��K�����M��uO�L+�߇���Q�g�:)�(؏�+�>��/1m#)J�t-����iTe�˜:�eӉ����/��Aƹ5��ùF��}�Ug7Q3�z�+ݿ�}1�8�<O^��C[�w�je9��A�y<Z#I�Wr<pTe��B���i҂�ʵ�"�UӖjyZ9���yZʄ������gh1{��{aO��R<ER�c�۶�~�:�����2`+�}����]��HG�Y���ݩu���}Y}&IO��*+{�޸�UbX��x6D�V�ez��"�-�$U��u�0l���l�̛u8���)r�Zس��"j�E� �a�O-����q>�T9�w�>?��@����LL�q���%2��n?��E�FF�a�͋�[�VE@����O�'w0X��KP�0���I�1ο���G����z�I_aծ�����"��2V���g	<K�#þ���޻�|<�ỏ��}�"FV*|�]WT�V�����t=�d+A�O�i�:���$�rƪ��H�=8��h
�����teV�j��pE��fz\�Խ�n��3/0�w�J"��غW4��~�B�eӊ���f"
�����V��p��Ɛ���H�B�#�P��[��>7�����t��x��m;��ن2�ޖ� u/��KBp�)P��,��B{A��5��醑�~��ݛ�oͤ2~$�˸����W2����-��9�cRGö�����@�Zy�~����������'�Ӧd6_#3��ϗ�^o��	Y��=o[�ެ��q�;b��tQ�_��Ɖ}�+��DP���U��	���^M��PСZ2<�k[)��؅'�Y�G�1m�	�y��q*�_zu�=E�N���o���A_\P�1��3e)���=��N�^�.��r>(){~w����`k���ȮJ�YxJjWR�i.���I�f���f��'��VwYs�:ShT]c�;?W��g������������x���`����O��U"v>��`��wr�S�&r �L(��T��f)�o�}��޻5s��/,X|�Yi�(x3�+�JFfωA��S"�}�;r%�g�?]�Hq�Al�hĤ����tjv�q|�P�{�g7/�Ko�,�<e-t{��{$�y��5�����틳�%�YԎ����=mc�ޢ8�#I&�"��?K5�E}dB7<W��C�*����Z�8[��v�3nV�B,���&�Ϥ^�s���ik��*�H��ў���L���+��|#�e`��k$}�}�Ӭ��ìŶ�$J�?r�}iɅ�*��5���������3���_ƈN�\J�]�f�ef�V�P˭��G��`nE�~%DmQ��P8r����ݿO�����$=Z�o�N�MҢ�Q��s�
��^��V��3�_��~NIs�1*�zj>��jى7�W7!�ui�ݘm(�|2����� B�i�[��s��m=����t:F�߫B��⛤��c��L��T3T�ϫ����R�v)m���?���� Ga��f��H׾��ʭ�)��rk�)J�^o�f��:�F�n�	�H���Ӗ�����ػ�Z6�,la_b�D!��ɑ�5Ы��4o��jHGL�*O�0�����S]������>�~��J��+��"��w�Bg���WS-R�Q�0;gY
�P�O�ܻ�Iyz�ZD�z�aQ�����2k֮(��H�=$������Y��p��@�*���/�ػ�v����"{ƾlj�P0������x0iD� ��e*JW�� ���*eZ������ �v��74�ʟ�Q����N��F��g��p���9�<�ߤ��a�ؙ��Q�!���d������C��CC�$ۼ<cb��V%w��y��yK����u��)�Fuǅ ��O�N�n鿅�r��J$��y�Rՙ/���w$]�	���T�%���Q�߂3�+��s����Sz7]���0ePJ��7ir�0a^�Z�{�!�tE`N�5�+���z�@}�I
����5Ǐ�RW�������V7M�����=�Nh-�dİ�_�(N�Z�E}%|L;�
�h��g
�u�GDV��y@�P�v"�7O��9�~0Q�J���N�h�ӴM�B�8��ۖKU2l�~�n?����\xդ"@h
ކ+D����Xh����[.�=��W�7���r��|#��ja
���6������Y=,��4���;i�?�<�w�\��"Mr�s9�Si,"���v��{�M��Il�\o�S�!�N@z��� �V#���/����qj�d�B7�=n�+���극@7t���������;9	���$���(���M���a%�ۨ��Fs�5}���b��4p@8�5 �����귫І���_b�ث}Pm1���]	�0)︪H��׆��?i�D#�Ǘ�
Q��Y0h<�y��Y�)�SQ^` �����-�Gz��pʺ~�$��6Sw�l���1$ +��zE�eN��b�5��mjA3��f[BL�Kw�F7�*jU ����[ډ0U�-�"0�n�B'�ƣf���=�N	́�Y����D�I1�������:������nN��IZl��N
�?�>��Td)� ��/�*;�"��ͫciA��SlՀ����ی��U�*����*MdM�h�� ����7jh��]S���=�ws��+,�3���/�H�N���&��p��p���ti���
��¿|8���f���@�0���>N�
��O��JC�����8�G#fT~��*�	�C�4?�� m�A;�[�)�_F0n�h�!AT�m^��` �t���r'c��I-��2���?~W�jOi��l+ G���J�ݙ�la�m����p�Aİ��j14{�����,͒`�5�~n"���_��i�����1�,J
��6kp��k�_a|O��S7(�N��h�	��BW�������3�z�L;���q�hq1��)�Т��@ZQ�����Y��0��W��ldG�D�A|��5G�]F6Z�?�f�o��t��2c��>U5��>����_��9�-���%)i+�X�OG�O�Z�P��D'��T"��g�����TxM�b8���٨�*��F�<y�hl�.�-�#�9�J����w���_E|III�}�ity���2��T"rJJe---�����/>8��dvS��"-�(�1�iVI����k54��uQ���)Z�s�5���
�;����l��O�����B�0�.�
�z"�0<�Dl�p������y��F�]�wп�����x�Ȓ�4��d��5��q����P��8���`���0�b\Rol���=?+a���X҅ �u(�F?���8�����_
��bV��j���C�9�]E��{j�8�r�q8���GԴ�������W��;���2f:����;��h��ќ����;UQ��<^�����y���4V��#w�!ײ��2��8�,�����G�T۸;)[���	��ꨈ��ƶG�?*"B�2����֢'�Ջ��v�a����Ш3�Z��|�*��������x���S�V���&Ԋɢ�K�����+��F�bX
1�cc:~P�Ѥ�o_�l�v�&d_����^��^��E��PWJ���+�C��Ȑ�!���1����ii����)��B����Y��ֶ����_d0��B�F�0)֘�J�_�5�9�)�
������`p��7�t.��{{U.\ �p�f����H��U�(��G�����*��D)]Y�sz�B��6��[�w~>��ŋ��W�����yP�1��P����+��i�9�Jî���n�8��{.4E��P�ɷ-��>x\`o��j��~��=�N�� B>&8��"@�J~���_�=�I�2-_nn���V�R��Q�`|�x3�eg{�o�"g`p�3��,O�cU�qS��a&�(��P�D^����^��~�ҫ3�L�0���ٙjM�����R��^�I�|��blwW^���������/�x+�\>�z[̵��!��i;���C��Z�B�$��ح>'ҕ2�Mb�k�c�ga��ԙO���5����+X��D�m��}�h��`�Ì�f�M8[a[娠8/
��)�@���q��&��L(��q��(����maj�/=g��V�����Ԣ�s��^���Ȍ��S����_#"Z��#�AĮ� ������?�~}-+h�ͬ��{Tm��,�8[-$$�z��o����в�c�A��!׸}�5fuC�T���O����m��33<��LN�N�s��=��1�� ��#�������p�Y�߳��1�@u��?�d�N���ER�d�睡��s����E�]ǽ7;��ݼ"�/84�����Ν���Ȁ��L.�ɋ�Q��n14Q�v􉍻���ލ+�i�����FY�y�7������w�{�'��ee�g"Us�֚�����[��B�Y_��K���-�p}��]���JIg]��%<��o̊R;gM���4�^*]��s��i���]����W7�p������h�a��j��=s	Q�шg��ޫ�9T�,��b���8}�[T/��$i|T���VIi	��k|w���Z#�M�&Y*���boo$6J:���;7??2""��˩fܑ?I�a:F!;����ffV�+�L��J`}v���]~���!T��]9�T�	ɢRfFƋ���222&\��Ŵe66>�׫�l�lni�`+G�^��f��i�fuS��cbf��eP�(���������ˡq���9�ȱ�Rq˗�H1��o>�����;+��(�x��"�˃[�𸘘�����TTQ����9�rv�k����=7~1nw��2-�t�f�Д����V9����{e�{ص����h�U�2���bhi�i�X�SpgmQ�m�^AᶒV�%+����ohߡ�@��h���z-�3����O�4%'|�'�{c	�$�!��%��-��.��jVP2]y�o���z���@|Lɻ��X�{ff&q3�*�'�J��X���)�U،"�R�Z����������!��T���d�9r� ���7�����(�H�(UQ���g����v]�qq9�B�����eB�-��y���Ř�_r�/�<9�Ⱦf���z�5�����l����/ �ٳ`��@N�q�q���y�{{.y��9 ߽,����Y�V&�_!:�C���x���t%�Ɔ�L�O��fr��ӭQ;�=�noo��`_�{�����$~�+��"(��5�����W�%�����kS�D����۸a�U@E7�����Ł�+;8S{-{t�Q�Q��ji�|)����P4>�i�?��#�z\� ���d���gfeU��K���,��Cxt���~�vj��IQ�kjh�KAЛ���a�gw�b�V��A�
X0��
S�A�sǰz˃ѡcZ��c
�wl*
�E,rd?T�M�Ё()y���1Y�'W��o�f�T��9�����働t^bb�
/�����
����ڕ��^-� R�4����"$��v,@������x���Y�������Ƈ���Kf��K訠?�`�qe2a(����uQ��4-���W��~��������Cu�o�4*6����,���"��J����-<��Ty�p�r�+墬������BL�/W�*�K1
���=�<�?2�#ޫ�l+Y��t���>{D�/6��%ך
��zV�(?�t��#e�!�B�u�L�5h!�3$�l[�{h]� sM�$el#w��m������4Z���Z����T�0} Y�.��qk������ }��	~P�L1�<AI�uwafc����J?8�P!�=tH�Z'��MC���TUY��>�J����\�2Īƨ��D�	h�_�E~H�
z��ݯ_��dq7T�Օg�>�^@B�룅����?P�ػ�� �����K�?��&��0pY��a@u���,����{�/��Z/�B��>L�mֵ��v�]�.����984����V�B4#�m6�i*�ÔO�p���%�����(Z��$%巶���E��v\������%};I������Dj&}^ ෶X'��+W���vě�<��(����S���L��~��{��1�ˮ�e��W<����dA�*��vrDC�
7|~�� �%�ٽg�_��޷wM�?���/]}u\T]-"�tw�4�H
�)CI*�]"JI�P"%  ��"�tww��w��}����7p�9{?�zֳ�>w��z�u�?g�h�mk~���d�H"Gr�T�?S�YPk�uZ���&����X#Z�av�ve���"����Xw��d�^�:�uu�t��k>̄��
�U��%g�����v_
����]p !f��ى����2��_�?���\��|x.�S�(4=]�C���=���>�%<�
�U(��G?:݁)m*7������vz����|��Eod����2�iXe�#��Zq{ϸ*ٽHHmS�J���N-p�����ЌmM��w:�<��xRE<�|N��j�/�%������U`��*��C(mPߑ_�=���nҶ�����Z�_�!ۄ�/}�"�S	D1	���0��-�B�l�}�at��;�5�J���T�2����QfK�w�C�r��?��}p��g�%�:n��o���h>}���ͽ�X2�Ϛ�j--Mz���f���7�~���r��=��I�583	�Δy�Ejzmgn��Ћ,����|<���Ζp܁��Щ������R�|O��n�f��&�N��n΄k�l�aj�'6h��A��4>"�J�%"#���S�A,r�7��/鴺-y\�''�w�oT��~��E���޾ɼ<�_�?W���!*����/O��%C97y��7|���K����k�~L�҅(e�8m��i���M����r��-�[Ai�$6��k�?]W+M��L���8�/�så=��n}����,u����|��W����E����p�W�i��??Q�/�T6#(��h�ْ�R�JG�;-�����5\�e��ؚHJ���}�7�>V8��!)NlDa�9���3C:�ή�>�/�� � r�@���$�&l�G�ՙTooo�p�ZoW�:C�m��i{�HL�k iw��^b�1o�c�Z
�?��x���92��=U���x����c���P�l�V�tdA��ȝ�$��r�{Mjx����6IQ9�WuurR��~��>������}�S
��`t���!�Hp���A���X��6a���d��H�7�Y�
���$b��y+�����j��D���)��+YLo�Y)!��g����D2w����Q�BF[����/V������t���VO�f��#"���}����8A�T��g�U����#.m�郱�>��@���57��j���Wlͭ�.�6��k�j��ք���o�b�P�Dغi��_�����뀋��J�`�
��*4�N��ъ�:`;o.3R��{�6�Fe���lw�Σ=)�H��1q�yW,���
[�X蠺�+����N���xW�b*��y���h��z�pi����ﺝ�AI�ǳͳԴB'����Mn���n��fx�2U��F�d��I_���Zhq�����*:�#Q4���.パ1�ݭѐ�LQ��)ܜJ���]_�5T��@ 4e�ld	�{���@�?�}I�ؘ��G8ˀ��R������_�� ©���f����h�4�ݓm�����rt���>F�)g�^ (A�BSx �Z��1'��?���ĲM�f��<��VDP�����9��G���?�%)k��r�{�g�(�x�ZS�pKĂ��sC���_�X`�C���ۜ_8��P{���mx�Z&�"�{_�O��5TM����\�`�
�8z^�W��x�0�����l+vrr������b<5�It۪������.��;�}��Z��v�o�\�e���Y[�~+��AXDt~|��fBt�8P�D�6ik�8��<�v�K Vq��T�^�9�z�V��|L��{���d�g�'̿�KtYQ�l��J*�a���ޮ� a��8E�^�B��3 @�� �	�����;L���G��c������gi(���MX�������AT�56�F?qX�z���A��<��%`�3B-y�ż�Q������j��:L���擇:��9�~��z�}�h�ZU���eL=U�{���.��Ff�f��gv���9�6��e:���foD\����CB��f|�N���*���=(O�!�~�>e�c��xQgsp�-Qٓ+,��ǳ|(&�OQR�O��G�ύ���r�q���9)))�' �ń������Y�=��'�:�APf�MBm�P:f���dS*>���6��嶯#��{&��l�L��D�啕� %�+���>�m�:��� ����Ὁ�Y���2s��������VM��Bv�;��Х��"%eeK�7��BAGB�5�	�f..�����L�Ԓ�Nu��u�^�4��gW�������������P̜޲!��Tz�}�ob��+��u�,��9�����:�}dF���g0aL�i��%֬X�ٟ�o�<Bղ��
�����I@F�y^fK�H�, )�V��Pqھ��a�V����-q�Q3�W�m��r)��%=�����#7\K +��94-� !�Jfhm��V4K�����4����'<��C:�m
���B4�J��X]��IJ��/U牚;�kc�d �̒r��X���Ub��̍�i�e�����*�'������F7L��&!��+.�p�yi�= ;$uSY�y�G�*=;j�b���$����2�(�́(�ql�)�����z����L@ 1�ݛ���)G_�����`��~2,�~�S��r��������mB�e�fl�|���Y��MW������fNŌ�2����V��sC��Ĝ��~\1bI�y���C��\��)�"Z%b�F��;oWc�g��#���t*�,�͕D:�H����G�yĮD��W�A�`&ϨO�z��#S�#�������\����W�� �lw����us�_�g����H��i23���9�П���!F�V޿�^��Ʈ����{/�Im��{ҹ�Cs��a�Gv��mZl�7�c5��3Ep�ZdogA��m!����ek�#*B��6|V����Nc��;�ĝ:A�+Zs�Y��p�Ą��	�<`��bdddM[e����m�>��94��T�U�z1��������_�G��x>{~Hʥ��WJ}�;`@iy����~���Ӣ�d����w~����o��X���,p�X���z�IAX���p�痣�?|/ҁq���d��������(��TL�[Ș�`i�6��u��ׇ�V���pݸR�4,��&���a�H!n��ͧp;
�>��2�*��׌

�4�Y�fJ֜�C#_v��Ơ��T�� Q!щm���î�m�*�U��J�-Xs+X��W��ٔ�=�T�4d�Gވ�k�P�Dޒ����(�Gv�=$*Q��tnr?��y�L���dɭ��v��]���k��s��x���׌��l��\C�^�	B��!��d`KPP�N� tXNe�[��M��������}�S�>�|1R�dlt4��w�ߗ�I�ϩp~*{o���Q:�<}|ȳn ��g!c�U}3ө¦&����P;f�ϳ�Hv��6�����A�`�2�3s����^FO�l��}E �6L�~傇������K�~�Sz���1M9$���8� y4��k��Bww���o���ȉ���?�U �[��t��G���e]�2#p�x����S�m<!�	��� �4��'tE�����kmV��;��Q�u`ya3ܝǵY����^�ٱg�lOT��/h/|�<�%��%x1�EQ��N�"a���YU�k͟lt���<��y�`+�c�ː��T�k�����|���USe������	]z�$>4�hfI���"	�W;�"�_����	��Q�j�cD5��������CQ����:b[�r6��r��M�1pw�!���l�a�����[����<�i�� ?V���������[(b8��f]�^�w-���&���Z����3|u��]�WT�����ʈf"%�W9�.t�\i��Ũ��y����oN֗��n�~X_���|ck�������h	�KZ�ռ�n��166P���r�+e9HZ�������:���ubf��?}�MO��3�z#��ж�	%����������
Њ�����e��?��5�O���6��|����#��Xr��EMC���W�7P��5���{"BCS����?)qʮ�$����Z\��@M�@-�����{vE3��gf�gϚ��/��pj*m��\o��K��e�D��i�'�����v��_(;�Ó�׏� ���-T��wQ������>  ]��8���2��nK���Z#Q }�(r��%��rJ��)��|�V�}��	��ѥ��ez;�mS����ώ��w{_�)�7n"����2���j5�sIh��ɯ�|�P�ܕvv�+Y��	���^�����a��Ә�ز<���g�x��SP���́�w4���c��sIa�ج�� -~��*�c�G�Â�Bo����{\&l�ؖ�੝�������V�����]͈�����'n��D��	�ͱ_�""��`���D,�1yr���*>Ni��l�Bڎ�D!�T��05��5�k5/,�Q,����6��D�S@����Q�K\n�p7wq�?dkFpD��ar��4Bd.�P	u������HL��<�T_߀�y&�͑4.�˟�-���ߙ<7ܖL`�滢���Ox��J?xV�HH ;п)è`��{���w��4�+Ft�4(D]����V�wVj��*  ����Ն�'��a-��yԛ�[�#a;;;��� mW	/'��:�� �Ŝk�j(�����d1=:�d�ܷ�[�03$�f�j&��C���3���8^�ޞ�8��ެ���`v\�UM���卽ۓ���pD�~l��g�su瀞4P_W��::fJ(-'�E�F�A�]�/�)����=�������ӝ)<�77�5���iH"u�?�4/8�SΝcd^��� ��uA�q�|s<պ�-��j]dx��ٳ��Uk|���5��d��mҰ�����>0�
�P(l���eb��٬�2���`>a�Ƃ�6qp��R�|T�VHt9���?\gMg���g@�kS�}��|p�G*N.uX�I�H�����Bwq���Kt�a��s^*��*�2
q�Iq)��j���N�$�켼�u�����j��ݽ���=�e����?�~�\b����iļ_%Y���{�y����=A�@dd�s������޴cM�c�h/��H}}}�ggc�������]�����r}����?ha�ꝡq���] ^��a��ެ������5P�ΰC�`�'�@U	t��X�7D��D�Z���~��.fNT"<ѓ�!�@�s���UW}��[9g)�uǺ�r22�����C��C=�zEv��ʽѥN�f���2j��L�� ��o}��g&wu��ֲ�Jo�d�=<�<	e�|)v��ZD�yD{�9"m�
#+��\�r�ϸ�w�
Et����1S6ZT���ڣ����͓�4��DG�R�z*�	D�m�=S�p�%�L3�~��Z�9���)n�< �*�[�T�)�[!����l�ht�>�H����rd�y�&���>A�ޒ�X$@�@%w�zAK�%�h�a���������s4�ڜnh}y	i���/����G��^�]��X��/����2�KV}��8-���Y�RlkYsӪ;2��<����L���Mq�ڿ?������|��t=yX�ˣ�L�7��]&۬�5�Y��5Ȗ����ܸc�ͤ�.����2%$�P�Vi�)f!m�ޚ��~M3�{�1-��ά5�#�]r^#��������D��`�J�X�y�N���A���آVc���qR��8
��c:�Z�P��i������H�9P���>�w�U�Z��_~�}�ts��\DWRj��n�����^2�2���*����4g;��GUp�zw�ߙ1m��}=��ĸx \z=Ǣ������c{ȟާJ�׆���E�*��@C�	����$P/��Bk٤��nkL�4�x��z��q��_������GP< DJ���i#n�i�
����k9���襳?�6�y �"��ōԦ����YN�h%��#�������0�^�_BS�\k�m�6im�("CaҠaa+�,"��	�2�T�,�BS�0�kg�c�
W\$蓙0-��?���;Wnޛ�9}�i��3�'r��uQw����"�\��d4���(�t�D�X݀� ���$9Z,@��&a�0��Hqcr�wE��1@����\�����%j�%b�S���`��%S$-�
���nc��F�}�ހ�ڢ�7h�H'���TY 0�I��N��0ǩ�yq���Ah^��R�5��*�^�:W�IN4,T���!1��}��Lz������E
��
C�R�L��@a������3�³��Z���b[�sO �(i����Bomd���C����9�9e��C��8�k!�W�]̶���K����H����)���ې��BxcU��l���Z\E����
���Mx
s��<b�(�'Q���:�O�c�S�_vH�3;�Q�jA.م�czc>�ﺳx�G�S��V�eAM;eSkQճ���N�"�0U��6ʬ����t�RGE���n�@���8���d�k�eZ"3�����ŝ�{Pf�z#7*��T]�Rf5���
�N�Yd�TzuX��
V�y8�F�.��w�dК��{dkHttt�����j���݀�b�'XX�s1�d�����0��54�It���TהԪ�	��f���g���S�R�ܣ�,�i��+i\����I���ճt�EPÅ?u'���*���ʖ����u�v��ߺL�i�Ԅ�O��ќr��gN�ecv�*�
n$���xR�Y�dr�>�_�"���d�\WMT�J,���i��|��K�·h�Y�c�w��z�	-�z��wM����ch� �k=�g��~"/V$�=��/N;P�E��|�R��tG,�N�@U�X��u{#_��E%�5:sQ���6+].��cU�
vA� �a7>fm���n��~�B����]ה.�!�y��w��w"fMC@��Z|��M�1��޲)�T�����H�1���Oi�g����r*�6��'�O�M�Jw]&�~,��˿h�zΥ�mE�Cz"�B$��������Mn�"��?Mi�â=c�J�fҬ_�n*�p���� `|�jNX��Gv{�摙$q-w����h�[����f��2\L�q�]!%��r1�:�U%� 밧����ˤ(͜P�������w
��s�dz��zf���O�����4VKq3�b-V�N��hߣ,�B�UH,��6i�>`��ט�sL�z!V�RgW���m,M,c
U2|-E�����	�1U�$!U�sŗ�tr�KwK�+�6�Ϸ���ې�cdF'�G��O[$MwiOȫ̬ʴLC�ph���t{"W�""BAy?��^����E/샳%�B�6��=<�	N�=O-�CtJcȉI�+P�n{�{�V��^SI��.��֍3��m�U+"���,5�	N�98o;ɯ,������#��U]��k�h:�2�Vr���^�uO����*�T�R��ˏ_��M� ����\Dzo��E�U�p7jѢ�D�Y�B�g����^��D�J��fO�u����]{"�a�ܴB�~H���MH��jI��뤣آN��4Us�b�f��`��9?4������W��m��4ʇz"�2�����bi�
U5t�9>_��*�b�&h�W��nzR.�:�4D���?F�!�ԛ�V��yo��ĵ/1��$}B����<o�}|�m��:�
�t�Ħ�mJ���b*��O�|��Ut,n�#�?Y���	�L�ɯG&�9�YM~��6�cv�@�B�����z���� ��f�c{��m��Ͷ��170�j�}�OD��O��o\�MplmS�.�勬�o���P6��'{yox�{������(��Z�.�u�z�s?Qd��TW[�N�������p�Bp�q�W��Tv�H/�m�����D22�9ѵ����&Q�X�mBoFs�X��*J ��^I�23ۀ���P��8�z%&��@�\�o���]�_� x�&��G���i�����J6*�w!���1���ә>R�޼mbK��:m�]>�Ҍ^4��:_#	��tC.�����P�db%�*��5���ǥ�`%��B�7�����c�ۯ�̭_?Q�]ŗR� ]���xP����B�߫z"�ˬ"mL����~T�MwII\����9�n^���?F��� ��ݙ�o1�VN�V�6>�B��m��������&�3'5��k�i�왕���4)vmH�
3)���Z�5�g�F�2���+)�+�Ӊ|�3�o8e�Z-�3p���s6J�#&�z�ٖ�B>f�֏�u��gI>fI�SS� ��u&�(�N���s��M��|{�	��HW��_����a�<��0�>w)F)�g��B5�xw|�&�������M�rV:�~O�iv̜�N�;��I	�(E��bTp��p_=��z�iJ���]lؑ��޳�V7�k�����{��#��� '�mJ���F��`�`1؃ׇ7ח���R:��;v�Z�Ab4k�=��6�3�w�~"�L���/�y�f67���ÂB�+&9���{S9�B��{]+3bq��1B�xC�ߏ�cx�˺�ٺ���X
t�
�ܺ��uJJ��L���QyQ�mr.W�*\9��}2��(2�n�w��ݙ
��vcG�_7ڑʿ���D��̢X�U�+I�����_��S�|9�Nd�3J���
~����Z����� a*�$����[(�����$],�~:ř��~|rِ@��O�%Il%�����C�EJ&��B���NBx�)�VS]�DKi~��c(m~�� �Ĉ�9q+'b�$'��ن�-`�	�����d����yS�ǚ�S@�ʽ��c=}S,PB(�5&�^]��1v�_u&���dd�I�i���Ӻ·$!�d�.�q�.�j.���,ۨ�d�U��C�Q��?�q3�Zo`r�0��/�����|��)M��t\��B�c$�.Q.ͦ�d�6i�z|r��<��-څ�-j�~�fe�VUxs�S{B]c�����������\�G��#�1���3�����H#���7F+�=�Lʲ�jl��/�572��\�.7�N������!�ZD[[�?Jw%�'_�!��)0)���>Sb�䎒bJ�����)O&�I�
��c�WrG���,�i^Jh1C�I(�bQ7!�|�F��Z�*h��5��n�����}���w
6K�����s��i�@�'�߽�_�\����'�DQ��D�K�I�JD�xI�<�~4�F��=�7O֑��l{�B�PO;;vdD�,���5�%(v�HapL�M�8�Z��\�}������!����xy<M�R������a�������"*
	X�оNLN~B{��x%��Ww��7pt��(���8
��(`���	��y!7����{�O�~��ǋD��K���멽���$Sin���]��Ck͇�cJ�6� L���rA��c,т}Q�9;�����2�\��t�+���?1��e7/'�����fTr�1����tJ����iE���8�{f���v�]1���c�5��9�)��"\��GıL�'�m������]�M��d�w���{�nO�I�p���d>�������:r�f��1���քK�Nn�ԉ�)�UCib�����,�/��1�Bsw\뉬��%�$AX�V!���cʗa��| �Q�ѯ�!��/)���W|�����L��� ]��w�uO��yWz#�Ƚ����v��VF̊�N��� Z����G�y�X ����g�lX�&O�HR�:p:�ݻ@���O�R�e>rj��)��?���G������*��"��h7�>���R􊨷��/�~��d�UЯ��D��B�Vx�@�G�ٝ��
�@.��]���Lv�Dl��{,,�%������G�!�B�~+I�`���S�wg���uvٸ*������ڃ��9m�he�wL����O'�N��HT�A��8��죞�{�!t�������!k4n9?���,���Z3�À�_�}Ԝ��U��o�?�H�!��$���x��-m��A?�"�ݟ�+ʪɔJ���PK   ��dXl�>��  |c     jsons/user_defined.json�\[oG��+�^�=�KU_�&K�F{lːl#�"X̥'&M*� �߷zH�����G1�r���U_�7u���l�۝?{v����4�]�|s6?��7����~�^��~W��ޟ=����xS~
{�iv��z���5}�.�����7����E�Y���v�^.���yty�y֖�{??[ЏgR5W� rf�׬�b�R�A �����fq��/����EM�nA6�c�Tm�F8f�1��}��w�����_� ����Y�y�l�Z�/���U�>{���j��rq�,�X/��Z]�����7�_�����,�V�_v���Us��,��_X�/��_/��P�炇_,��W��������v�#j�e�÷޿y����y\�苅���r��o^�+�b1K썿��A��/Vg�U��0(�RM�T��}�6K�_�?,����P�*y���ِP�*����A��/s�����7+����rXhߨd����a�}��y��B�%�T������9>�|T��ūa���b/χ�FlJ�=O9@�7+!�䦌U�K�<��"�\}��+v�d$ha��a�����s��	Z&S���Y6S��ڷ��k�H5�R�6&E�T=,�ob]0ȑ:�ed$n�L��QFdJ6/	]�)uغT$v�L��ƥ"��dJ%���Kc��k�_J�����T~�`�Zi�J��"0P�e����U+K^7J���n�����P:���B)�����V��(�����Ur���=$�׿^�.֟8���j�|����v	t�g�\�ڲ��6T��@��o M��'�_m?<�S�X�T��_��N�/K�q����?��qƋ�[��_of�~��>c��ZO�X ��T�"�j�F]�F�3���o!����*�*4�A�Y��ٖ��H�R�P�8-��w�p����9��ϭ.��.�'ʫj+#H����C��U��K!�#���F����J8���	"�TR�<R}q����IÑ=�:
�ҖO�Ű����R�BHp8	b��G2JC1_��߼�"�R��
QX�4��eR)'��I��r �V�qN����P�)y$��D�$53��`� ��ԺB��\U���5ЋW	�"e��� >!Q��\ӣp�17D�����v{��)b�Ai����h�H����w���u����|�}C�PV@k�i��f�aP4��\�=I��<bds�6�H�Ia�����I�"�f�A.Q�s%Ӂ<ɿ`ds%�\Eb9�Bs w�͕Js���!�ϕJsշ�#F6W*�U$�s.+�r�dA��HD�@��	lA��H@?�d�i�"�P
t\�|�0IW���@&*&銔�' �ta:��Dt���D;�..B�`��ꂥ:�*�y�XG��$�DUE�wܼ�eJ��H
o�A:�^SP�?b�@{	.�ܰ4Jk����k���a���#�P.*�$��H���S�ث�$��S��}��X����
Īt!!"kѡV-G��o/��l%��A1����r���ql���?�*8��:b�Gױf�M�)�"�D��J���$� �N��^Ĩg�#��"�j�XHc(#�.��-=��Ż��w?0�a�m �.��C�U��X�}Ez�G,+t!�^�k+�䑆��	(��b�(>��s�T�G(�@U4b�=�Q����	��@�&�Ô�c��W������࠺"k씒��DJ� ����U�$q"rZu�������BQN�M�K=�[}��aP����
	��.�#������
B�c���J�U}�APen�"�a�t��O r�"�a�t�����9m'%D龙w$v�D�����@d%SDE|���଄H���ZM J�������D�Q��U�tV�	D�Q��A��1��x��Ho��MOe"�=+�í	D�O&���#L�}.A������4�K����]w��dS,EZz�b���)�"�#B.K6�R��� ��dR4E����z�ϓI�)�O r�2)�"=�4U<v���Q6R�wR�	
�D�H-�K�Ne#e�B]P��ML���;.�Da��H�~�K�����J&�kB��X�.@he'<H���\� ET�e�d8/��J��6b��QfQ���E��"��TN�"�m��!K�%*����U� �!��TN�"�}�KT*'w�ґ3'�r�Q�9� !P�	�f���u�@d�)�"��-@�,*����uw�	�OT*'w�[5G�\�R9�~.�Q�$� �u[T�3J��Fߖ�r���W��m��M���*�D���s9�Kނ�}���pFv�L�K���}���։���#�u.��]�
ﻃp�2u�N�]�r��}�С�s��椙���]���g���攖c�_����0������P�$���E�cg������3q^��#��Ѐ'*��������s@hc������}=ёi�}�fj���=��ɐb?I3�g-D�*�΅�����������z��V�k��,�Q��������zyKƞ�d���:;�_�l-�Pb�b�`r*_)�`	��_�.�~ydҎ�9��+5	q%���!ơc9����!���E~::�ZV�k��a`k˜��!p�]S�p�`���b�z�]�ِ�1����n�MNYT�r��sXrf����dum�o��V�:˝�p�E��)%Z�Y�p�֥k��,%��)���i��m�پ}4T��΁�<�U�M�U���x�����s��灾������~d%J �$�c����~)�|a)�S���Ѕ��y��
�%8��S]���\����ښ9�d�����lj�v�[lgW�f����M�����kIG뚁/�Yz2�u�W)����B�[��}%�}3#;��t�l����4�.�1MY2�E�6�'�Rʷ.�\K[U���qY9�rV5�3��6ei[�>L�YkW��ȨQ��Vʶe�pԭ��vUƬ#i����q{Z|�Q��;D+Uvs*���KR_[���wi�݉��c�sI~�]=�
��@j9�(�0~c�y�!.���<�ɻw�N��G� W����h�)���@��0��rlb�x�A[r�V�Ge���]� "�4ۑ��JJ�)~`/ޜ���~ˮ&8�=�� ��O��'9R�_+�R��P��_�o�Ft T�M��:��FTh+w
��r]���*�l��7��8 �	���#>!�#�X��?kg& $,�s�/ڔ���gU�������ߑU]��YW��ɤ�ER�`������y��zJ��Ήޮ��-oƻ���k��e����I��Zo�pT��܌��&1��@J��"�D+Y�־4R;ʷ2���y<E��RN<�=7T�� �(҆w�����M�e��+@�u֍E��LoZ	������bPW��BmYٴm)*J@�C�*�FQ������bvu3���l����ސG�u����'�%��@�Zٚ5Zz�jt��5^6�,s�K`i�o�*R2�j���QL�U
��b �}����:���~�a��q�N���p�E�(eֻ�w��Ou�J�A�2�~�N<�� ���vm��ꭁj)4-�2TF��TU��M%J�RuU�����������������P�R����L�9k�J�ԚZ�m���,}���Ъ*��30������mk.M)��6I!B�k�t���V{�5)I��sss�ZB^5S[�BH*�EX
�~���Z��b���N�m��VC	TN6�V#3Ws��tIEx_��:GY?߿�!�%=D#���Y�5��X!�ڶa�S�����?�j������@����]��ߗ��L-�����0{��n���jQO�w�D����;4��a�l��d�ƩRy�]�*x#� z����Z3����n}N���D_��
�zBH3�UL�@b.�!Jq%���f�t�Jd��nRo�W���N>U�cͶ?��"��m �= <c��[���/�0�������%Z��sN3�HՒ7,��ng��J(n�p����q����]��g���n�{a�7+����ٻ�D�}�;4�9�*[Ǹ��Y/)�U�=ş[��(���B�j#YH6Xe�d�X{K�z�a��6��G���)�}D'ɮ,�9j[��n$���۔�tXpk�����R�Q1�ŏ' R�q�e�~���� ���0�f��@�_zТ� 8�n���SNE�ѣE�jG[��Ʈ9=龑����j&�к��>z�]{Uk޴��f���PK
   ��dXqC,&'  ��                  cirkitFile.jsonPK
   ��dX#d�y_  G� /             S'  images/0700f4b8-b576-4b42-8309-cd2fa5470453.pngPK
   ��dXWC��)�  � /             �G images/093f54e3-331f-4155-80d0-fca9fbcaa25c.pngPK
   �dX����(w  +�  /             u images/1485337c-0c33-4cbd-84c8-adffa1b45f33.pngPK
   �dX��@� �S /             � images/15a77ed7-bb2d-43f5-af73-2cbf4ea4040d.pngPK
   ��dX� ���� 
� /             ��
 images/38cb4f51-bc72-4d24-b782-e5d855ce8001.pngPK
   ��dX�Yҙ<  �<  /             =_ images/4c2bed1b-fdcd-48c8-974c-5402e9db5193.pngPK
   ��dXv��� f~ /             #� images/4d249bba-3190-4770-b321-fb8fc027a237.pngPK
   ��dX��_8
  3
  /             0� images/57489f55-55cc-4ea4-8258-f1cf3d9c722d.pngPK
   �dX�A�x�L  �M  /             �� images/6470d57f-e26a-480a-a2b1-cdb1a5d6cbca.pngPK
   ��dX����H   C   /             �� images/8e6e9996-4250-48fd-a42c-980e5b13088a.pngPK
   ��dX��) oj /             � images/9b962a8e-14b5-4317-8666-1954827ef6fe.pngPK
   ��dX`$} [ /             �E images/a8bb870d-02b9-45f0-bd60-404fdaa8f6ff.pngPK
   �dXs!��}  {�  /             Q� images/c17cd92d-b315-46a0-b1f2-cfcea726969d.pngPK
   ��dX$7h�!  �!  /             �A images/c6364832-c854-438f-b38b-75bf2a0cd33f.pngPK
   ��dX/yR�c  ^  /             �c images/d2af519c-c065-45b5-bffd-6bf239de2b90.pngPK
   ��dX�'k�  �  /             xr images/e8452abc-1b33-4025-a556-b46ce3c60df1.pngPK
   ��dX�+�s;  z;  /             Ɖ images/f3037bb0-f56a-43e4-a2ff-17056f7c669b.pngPK
   ��dXP��/�  ǽ  /             �� images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.pngPK
   ��dXl�>��  |c               �w jsons/user_defined.jsonPK        ܈   